magic
tech scmos
timestamp 1769293095
<< nwell >>
rect 3882 3711 4248 3855
rect 5047 3711 5413 3855
rect 6202 3711 6568 3855
rect 7395 3711 7761 3855
rect 3881 3696 4248 3711
rect 5046 3696 5413 3711
rect 6201 3696 6568 3711
rect 7394 3696 7761 3711
rect 3065 2507 3224 2873
rect 8218 2822 8233 2823
rect 4357 2686 4694 2775
rect 6416 2707 6753 2796
rect 4232 2631 4694 2686
rect 6291 2652 6753 2707
rect 3209 2506 3224 2507
rect 8218 2456 8376 2822
rect 8218 1976 8233 1977
rect 3064 1597 3223 1963
rect 8218 1610 8376 1976
rect 3208 1596 3223 1597
rect 3064 657 3223 1023
rect 4486 984 4948 1039
rect 4486 895 4823 984
rect 6535 956 6997 1011
rect 8217 972 8232 973
rect 6535 867 6872 956
rect 3208 656 3223 657
rect 8217 606 8376 972
rect 3889 -252 4256 -237
rect 5043 -251 5410 -236
rect 6194 -251 6561 -236
rect 7285 -251 7652 -236
rect 3889 -396 4255 -252
rect 5043 -395 5409 -251
rect 6194 -395 6560 -251
rect 7285 -395 7651 -251
<< ntransistor >>
rect 4259 2616 4261 2620
rect 4297 2616 4299 2620
rect 4324 2616 4326 2620
rect 4347 2616 4349 2620
rect 4370 2616 4372 2620
rect 4400 2606 4402 2612
rect 4425 2589 4427 2615
rect 4450 2595 4452 2615
rect 4460 2595 4462 2615
rect 4470 2595 4472 2615
rect 4480 2595 4482 2615
rect 4490 2595 4492 2615
rect 4500 2605 4502 2615
rect 4525 2515 4527 2615
rect 4535 2515 4537 2615
rect 4545 2515 4547 2615
rect 4555 2515 4557 2615
rect 4565 2515 4567 2615
rect 4575 2560 4577 2615
rect 6318 2637 6320 2641
rect 6356 2637 6358 2641
rect 6383 2637 6385 2641
rect 6406 2637 6408 2641
rect 6429 2637 6431 2641
rect 6459 2627 6461 2633
rect 6484 2610 6486 2636
rect 6509 2616 6511 2636
rect 6519 2616 6521 2636
rect 6529 2616 6531 2636
rect 6539 2616 6541 2636
rect 6549 2616 6551 2636
rect 6559 2626 6561 2636
rect 6584 2536 6586 2636
rect 6594 2536 6596 2636
rect 6604 2536 6606 2636
rect 6614 2536 6616 2636
rect 6624 2536 6626 2636
rect 6634 2581 6636 2636
rect 4603 1055 4605 1110
rect 4613 1055 4615 1155
rect 4623 1055 4625 1155
rect 4633 1055 4635 1155
rect 4643 1055 4645 1155
rect 4653 1055 4655 1155
rect 4678 1055 4680 1065
rect 4688 1055 4690 1075
rect 4698 1055 4700 1075
rect 4708 1055 4710 1075
rect 4718 1055 4720 1075
rect 4728 1055 4730 1075
rect 4753 1055 4755 1081
rect 4778 1058 4780 1064
rect 4808 1050 4810 1054
rect 4831 1050 4833 1054
rect 4854 1050 4856 1054
rect 4881 1050 4883 1054
rect 4919 1050 4921 1054
rect 6652 1027 6654 1082
rect 6662 1027 6664 1127
rect 6672 1027 6674 1127
rect 6682 1027 6684 1127
rect 6692 1027 6694 1127
rect 6702 1027 6704 1127
rect 6727 1027 6729 1037
rect 6737 1027 6739 1047
rect 6747 1027 6749 1047
rect 6757 1027 6759 1047
rect 6767 1027 6769 1047
rect 6777 1027 6779 1047
rect 6802 1027 6804 1053
rect 6827 1030 6829 1036
rect 6857 1022 6859 1026
rect 6880 1022 6882 1026
rect 6903 1022 6905 1026
rect 6930 1022 6932 1026
rect 6968 1022 6970 1026
<< ptransistor >>
rect 4259 2652 4261 2658
rect 4297 2652 4299 2658
rect 4324 2652 4326 2658
rect 4347 2652 4349 2658
rect 4370 2652 4372 2658
rect 4400 2637 4402 2651
rect 4425 2637 4427 2698
rect 4450 2637 4452 2707
rect 4460 2637 4462 2707
rect 4470 2637 4472 2707
rect 4480 2637 4482 2707
rect 4525 2637 4527 2737
rect 4535 2637 4537 2737
rect 4545 2637 4547 2737
rect 4555 2637 4557 2737
rect 4565 2637 4567 2737
rect 4575 2637 4577 2737
rect 4585 2637 4587 2737
rect 4595 2637 4597 2737
rect 4605 2637 4607 2737
rect 4615 2637 4617 2737
rect 4625 2637 4627 2737
rect 4635 2637 4637 2737
rect 4645 2637 4647 2737
rect 4655 2637 4657 2670
rect 6318 2673 6320 2679
rect 6356 2673 6358 2679
rect 6383 2673 6385 2679
rect 6406 2673 6408 2679
rect 6429 2673 6431 2679
rect 6459 2658 6461 2672
rect 6484 2658 6486 2719
rect 6509 2658 6511 2728
rect 6519 2658 6521 2728
rect 6529 2658 6531 2728
rect 6539 2658 6541 2728
rect 6584 2658 6586 2758
rect 6594 2658 6596 2758
rect 6604 2658 6606 2758
rect 6614 2658 6616 2758
rect 6624 2658 6626 2758
rect 6634 2658 6636 2758
rect 6644 2658 6646 2758
rect 6654 2658 6656 2758
rect 6664 2658 6666 2758
rect 6674 2658 6676 2758
rect 6684 2658 6686 2758
rect 6694 2658 6696 2758
rect 6704 2658 6706 2758
rect 6714 2658 6716 2691
rect 4523 1000 4525 1033
rect 4533 933 4535 1033
rect 4543 933 4545 1033
rect 4553 933 4555 1033
rect 4563 933 4565 1033
rect 4573 933 4575 1033
rect 4583 933 4585 1033
rect 4593 933 4595 1033
rect 4603 933 4605 1033
rect 4613 933 4615 1033
rect 4623 933 4625 1033
rect 4633 933 4635 1033
rect 4643 933 4645 1033
rect 4653 933 4655 1033
rect 4698 963 4700 1033
rect 4708 963 4710 1033
rect 4718 963 4720 1033
rect 4728 963 4730 1033
rect 4753 972 4755 1033
rect 4778 1019 4780 1033
rect 4808 1012 4810 1018
rect 4831 1012 4833 1018
rect 4854 1012 4856 1018
rect 4881 1012 4883 1018
rect 4919 1012 4921 1018
rect 6572 972 6574 1005
rect 6582 905 6584 1005
rect 6592 905 6594 1005
rect 6602 905 6604 1005
rect 6612 905 6614 1005
rect 6622 905 6624 1005
rect 6632 905 6634 1005
rect 6642 905 6644 1005
rect 6652 905 6654 1005
rect 6662 905 6664 1005
rect 6672 905 6674 1005
rect 6682 905 6684 1005
rect 6692 905 6694 1005
rect 6702 905 6704 1005
rect 6747 935 6749 1005
rect 6757 935 6759 1005
rect 6767 935 6769 1005
rect 6777 935 6779 1005
rect 6802 944 6804 1005
rect 6827 991 6829 1005
rect 6857 984 6859 990
rect 6880 984 6882 990
rect 6903 984 6905 990
rect 6930 984 6932 990
rect 6968 984 6970 990
<< ndiffusion >>
rect 3929 3467 4196 3570
rect 5094 3467 5361 3570
rect 6249 3467 6516 3570
rect 7442 3467 7709 3570
rect 3350 2554 3453 2821
rect 4257 2616 4259 2620
rect 4261 2616 4263 2620
rect 4295 2616 4297 2620
rect 4299 2616 4301 2620
rect 4322 2616 4324 2620
rect 4326 2616 4328 2620
rect 4345 2616 4347 2620
rect 4349 2616 4351 2620
rect 4368 2616 4370 2620
rect 4372 2616 4374 2620
rect 4398 2606 4400 2612
rect 4402 2606 4404 2612
rect 4423 2589 4425 2615
rect 4427 2589 4429 2615
rect 4448 2595 4450 2615
rect 4452 2595 4454 2615
rect 4458 2595 4460 2615
rect 4462 2595 4464 2615
rect 4468 2595 4470 2615
rect 4472 2595 4474 2615
rect 4478 2595 4480 2615
rect 4482 2595 4484 2615
rect 4488 2595 4490 2615
rect 4492 2595 4494 2615
rect 4498 2605 4500 2615
rect 4502 2605 4504 2615
rect 4523 2515 4525 2615
rect 4527 2515 4529 2615
rect 4533 2515 4535 2615
rect 4537 2515 4539 2615
rect 4543 2515 4545 2615
rect 4547 2515 4549 2615
rect 4553 2515 4555 2615
rect 4557 2515 4559 2615
rect 4563 2515 4565 2615
rect 4567 2515 4569 2615
rect 4573 2560 4575 2615
rect 4577 2560 4579 2615
rect 6316 2637 6318 2641
rect 6320 2637 6322 2641
rect 6354 2637 6356 2641
rect 6358 2637 6360 2641
rect 6381 2637 6383 2641
rect 6385 2637 6387 2641
rect 6404 2637 6406 2641
rect 6408 2637 6410 2641
rect 6427 2637 6429 2641
rect 6431 2637 6433 2641
rect 6457 2627 6459 2633
rect 6461 2627 6463 2633
rect 6482 2610 6484 2636
rect 6486 2610 6488 2636
rect 6507 2616 6509 2636
rect 6511 2616 6513 2636
rect 6517 2616 6519 2636
rect 6521 2616 6523 2636
rect 6527 2616 6529 2636
rect 6531 2616 6533 2636
rect 6537 2616 6539 2636
rect 6541 2616 6543 2636
rect 6547 2616 6549 2636
rect 6551 2616 6553 2636
rect 6557 2626 6559 2636
rect 6561 2626 6563 2636
rect 6582 2536 6584 2636
rect 6586 2536 6588 2636
rect 6592 2536 6594 2636
rect 6596 2536 6598 2636
rect 6602 2536 6604 2636
rect 6606 2536 6608 2636
rect 6612 2536 6614 2636
rect 6616 2536 6618 2636
rect 6622 2536 6624 2636
rect 6626 2536 6628 2636
rect 6632 2581 6634 2636
rect 6636 2581 6638 2636
rect 7989 2508 8092 2775
rect 3349 1644 3452 1911
rect 7989 1662 8092 1929
rect 4601 1055 4603 1110
rect 4605 1055 4607 1110
rect 4611 1055 4613 1155
rect 4615 1055 4617 1155
rect 4621 1055 4623 1155
rect 4625 1055 4627 1155
rect 4631 1055 4633 1155
rect 4635 1055 4637 1155
rect 4641 1055 4643 1155
rect 4645 1055 4647 1155
rect 4651 1055 4653 1155
rect 4655 1055 4657 1155
rect 4676 1055 4678 1065
rect 4680 1055 4682 1065
rect 4686 1055 4688 1075
rect 4690 1055 4692 1075
rect 4696 1055 4698 1075
rect 4700 1055 4702 1075
rect 4706 1055 4708 1075
rect 4710 1055 4712 1075
rect 4716 1055 4718 1075
rect 4720 1055 4722 1075
rect 4726 1055 4728 1075
rect 4730 1055 4732 1075
rect 4751 1055 4753 1081
rect 4755 1055 4757 1081
rect 4776 1058 4778 1064
rect 4780 1058 4782 1064
rect 3349 704 3452 971
rect 4806 1050 4808 1054
rect 4810 1050 4812 1054
rect 4829 1050 4831 1054
rect 4833 1050 4835 1054
rect 4852 1050 4854 1054
rect 4856 1050 4858 1054
rect 4879 1050 4881 1054
rect 4883 1050 4885 1054
rect 4917 1050 4919 1054
rect 4921 1050 4923 1054
rect 6650 1027 6652 1082
rect 6654 1027 6656 1082
rect 6660 1027 6662 1127
rect 6664 1027 6666 1127
rect 6670 1027 6672 1127
rect 6674 1027 6676 1127
rect 6680 1027 6682 1127
rect 6684 1027 6686 1127
rect 6690 1027 6692 1127
rect 6694 1027 6696 1127
rect 6700 1027 6702 1127
rect 6704 1027 6706 1127
rect 6725 1027 6727 1037
rect 6729 1027 6731 1037
rect 6735 1027 6737 1047
rect 6739 1027 6741 1047
rect 6745 1027 6747 1047
rect 6749 1027 6751 1047
rect 6755 1027 6757 1047
rect 6759 1027 6761 1047
rect 6765 1027 6767 1047
rect 6769 1027 6771 1047
rect 6775 1027 6777 1047
rect 6779 1027 6781 1047
rect 6800 1027 6802 1053
rect 6804 1027 6806 1053
rect 6825 1030 6827 1036
rect 6829 1030 6831 1036
rect 6855 1022 6857 1026
rect 6859 1022 6861 1026
rect 6878 1022 6880 1026
rect 6882 1022 6884 1026
rect 6901 1022 6903 1026
rect 6905 1022 6907 1026
rect 6928 1022 6930 1026
rect 6932 1022 6934 1026
rect 6966 1022 6968 1026
rect 6970 1022 6972 1026
rect 7988 658 8091 925
rect 3941 -111 4208 -8
rect 5095 -110 5362 -7
rect 6246 -110 6513 -7
rect 7337 -110 7604 -7
<< pdiffusion >>
rect 3927 3725 4196 3827
rect 5092 3725 5361 3827
rect 6247 3725 6516 3827
rect 7440 3725 7709 3827
rect 3093 2552 3195 2821
rect 4257 2653 4259 2658
rect 4252 2652 4259 2653
rect 4261 2653 4263 2658
rect 4261 2652 4268 2653
rect 4295 2653 4297 2658
rect 4290 2652 4297 2653
rect 4299 2653 4301 2658
rect 4299 2652 4306 2653
rect 4322 2653 4324 2658
rect 4317 2652 4324 2653
rect 4326 2653 4328 2658
rect 4326 2652 4333 2653
rect 4345 2653 4347 2658
rect 4340 2652 4347 2653
rect 4349 2653 4351 2658
rect 4349 2652 4356 2653
rect 4368 2653 4370 2658
rect 4363 2652 4370 2653
rect 4372 2653 4374 2658
rect 4372 2652 4379 2653
rect 4398 2637 4400 2651
rect 4402 2637 4404 2651
rect 4423 2637 4425 2698
rect 4427 2637 4429 2698
rect 4448 2637 4450 2707
rect 4452 2637 4454 2707
rect 4458 2637 4460 2707
rect 4462 2637 4464 2707
rect 4468 2637 4470 2707
rect 4472 2637 4474 2707
rect 4478 2637 4480 2707
rect 4482 2637 4484 2707
rect 4523 2637 4525 2737
rect 4527 2637 4529 2737
rect 4533 2637 4535 2737
rect 4537 2637 4539 2737
rect 4543 2637 4545 2737
rect 4547 2637 4549 2737
rect 4553 2637 4555 2737
rect 4557 2637 4559 2737
rect 4563 2637 4565 2737
rect 4567 2637 4569 2737
rect 4573 2637 4575 2737
rect 4577 2637 4579 2737
rect 4583 2637 4585 2737
rect 4587 2637 4589 2737
rect 4593 2637 4595 2737
rect 4597 2637 4599 2737
rect 4603 2637 4605 2737
rect 4607 2637 4609 2737
rect 4613 2637 4615 2737
rect 4617 2637 4619 2737
rect 4623 2637 4625 2737
rect 4627 2637 4629 2737
rect 4633 2637 4635 2737
rect 4637 2637 4639 2737
rect 4643 2637 4645 2737
rect 4647 2637 4649 2737
rect 4653 2637 4655 2670
rect 4657 2637 4659 2670
rect 6316 2674 6318 2679
rect 6311 2673 6318 2674
rect 6320 2674 6322 2679
rect 6320 2673 6327 2674
rect 6354 2674 6356 2679
rect 6349 2673 6356 2674
rect 6358 2674 6360 2679
rect 6358 2673 6365 2674
rect 6381 2674 6383 2679
rect 6376 2673 6383 2674
rect 6385 2674 6387 2679
rect 6385 2673 6392 2674
rect 6404 2674 6406 2679
rect 6399 2673 6406 2674
rect 6408 2674 6410 2679
rect 6408 2673 6415 2674
rect 6427 2674 6429 2679
rect 6422 2673 6429 2674
rect 6431 2674 6433 2679
rect 6431 2673 6438 2674
rect 6457 2658 6459 2672
rect 6461 2658 6463 2672
rect 6482 2658 6484 2719
rect 6486 2658 6488 2719
rect 6507 2658 6509 2728
rect 6511 2658 6513 2728
rect 6517 2658 6519 2728
rect 6521 2658 6523 2728
rect 6527 2658 6529 2728
rect 6531 2658 6533 2728
rect 6537 2658 6539 2728
rect 6541 2658 6543 2728
rect 6582 2658 6584 2758
rect 6586 2658 6588 2758
rect 6592 2658 6594 2758
rect 6596 2658 6598 2758
rect 6602 2658 6604 2758
rect 6606 2658 6608 2758
rect 6612 2658 6614 2758
rect 6616 2658 6618 2758
rect 6622 2658 6624 2758
rect 6626 2658 6628 2758
rect 6632 2658 6634 2758
rect 6636 2658 6638 2758
rect 6642 2658 6644 2758
rect 6646 2658 6648 2758
rect 6652 2658 6654 2758
rect 6656 2658 6658 2758
rect 6662 2658 6664 2758
rect 6666 2658 6668 2758
rect 6672 2658 6674 2758
rect 6676 2658 6678 2758
rect 6682 2658 6684 2758
rect 6686 2658 6688 2758
rect 6692 2658 6694 2758
rect 6696 2658 6698 2758
rect 6702 2658 6704 2758
rect 6706 2658 6708 2758
rect 6712 2658 6714 2691
rect 6716 2658 6718 2691
rect 8247 2508 8349 2777
rect 3092 1642 3194 1911
rect 8247 1662 8349 1931
rect 3092 702 3194 971
rect 4521 1000 4523 1033
rect 4525 1000 4527 1033
rect 4531 933 4533 1033
rect 4535 933 4537 1033
rect 4541 933 4543 1033
rect 4545 933 4547 1033
rect 4551 933 4553 1033
rect 4555 933 4557 1033
rect 4561 933 4563 1033
rect 4565 933 4567 1033
rect 4571 933 4573 1033
rect 4575 933 4577 1033
rect 4581 933 4583 1033
rect 4585 933 4587 1033
rect 4591 933 4593 1033
rect 4595 933 4597 1033
rect 4601 933 4603 1033
rect 4605 933 4607 1033
rect 4611 933 4613 1033
rect 4615 933 4617 1033
rect 4621 933 4623 1033
rect 4625 933 4627 1033
rect 4631 933 4633 1033
rect 4635 933 4637 1033
rect 4641 933 4643 1033
rect 4645 933 4647 1033
rect 4651 933 4653 1033
rect 4655 933 4657 1033
rect 4696 963 4698 1033
rect 4700 963 4702 1033
rect 4706 963 4708 1033
rect 4710 963 4712 1033
rect 4716 963 4718 1033
rect 4720 963 4722 1033
rect 4726 963 4728 1033
rect 4730 963 4732 1033
rect 4751 972 4753 1033
rect 4755 972 4757 1033
rect 4776 1019 4778 1033
rect 4780 1019 4782 1033
rect 4801 1017 4808 1018
rect 4806 1012 4808 1017
rect 4810 1017 4817 1018
rect 4810 1012 4812 1017
rect 4824 1017 4831 1018
rect 4829 1012 4831 1017
rect 4833 1017 4840 1018
rect 4833 1012 4835 1017
rect 4847 1017 4854 1018
rect 4852 1012 4854 1017
rect 4856 1017 4863 1018
rect 4856 1012 4858 1017
rect 4874 1017 4881 1018
rect 4879 1012 4881 1017
rect 4883 1017 4890 1018
rect 4883 1012 4885 1017
rect 4912 1017 4919 1018
rect 4917 1012 4919 1017
rect 4921 1017 4928 1018
rect 4921 1012 4923 1017
rect 6570 972 6572 1005
rect 6574 972 6576 1005
rect 6580 905 6582 1005
rect 6584 905 6586 1005
rect 6590 905 6592 1005
rect 6594 905 6596 1005
rect 6600 905 6602 1005
rect 6604 905 6606 1005
rect 6610 905 6612 1005
rect 6614 905 6616 1005
rect 6620 905 6622 1005
rect 6624 905 6626 1005
rect 6630 905 6632 1005
rect 6634 905 6636 1005
rect 6640 905 6642 1005
rect 6644 905 6646 1005
rect 6650 905 6652 1005
rect 6654 905 6656 1005
rect 6660 905 6662 1005
rect 6664 905 6666 1005
rect 6670 905 6672 1005
rect 6674 905 6676 1005
rect 6680 905 6682 1005
rect 6684 905 6686 1005
rect 6690 905 6692 1005
rect 6694 905 6696 1005
rect 6700 905 6702 1005
rect 6704 905 6706 1005
rect 6745 935 6747 1005
rect 6749 935 6751 1005
rect 6755 935 6757 1005
rect 6759 935 6761 1005
rect 6765 935 6767 1005
rect 6769 935 6771 1005
rect 6775 935 6777 1005
rect 6779 935 6781 1005
rect 6800 944 6802 1005
rect 6804 944 6806 1005
rect 6825 991 6827 1005
rect 6829 991 6831 1005
rect 6850 989 6857 990
rect 6855 984 6857 989
rect 6859 989 6866 990
rect 6859 984 6861 989
rect 6873 989 6880 990
rect 6878 984 6880 989
rect 6882 989 6889 990
rect 6882 984 6884 989
rect 6896 989 6903 990
rect 6901 984 6903 989
rect 6905 989 6912 990
rect 6905 984 6907 989
rect 6923 989 6930 990
rect 6928 984 6930 989
rect 6932 989 6939 990
rect 6932 984 6934 989
rect 6961 989 6968 990
rect 6966 984 6968 989
rect 6970 989 6977 990
rect 6970 984 6972 989
rect 8246 658 8348 927
rect 3941 -368 4210 -266
rect 5095 -367 5364 -265
rect 6246 -367 6515 -265
rect 7337 -367 7606 -265
<< ndcontact >>
rect 3913 3467 3929 3570
rect 4196 3467 4212 3570
rect 5078 3467 5094 3570
rect 5361 3467 5377 3570
rect 6233 3467 6249 3570
rect 6516 3467 6532 3570
rect 7426 3467 7442 3570
rect 7709 3467 7725 3570
rect 3350 2821 3453 2837
rect 3350 2538 3453 2554
rect 4252 2616 4257 2621
rect 4263 2616 4268 2621
rect 4290 2616 4295 2621
rect 4301 2616 4306 2621
rect 4317 2616 4322 2621
rect 4328 2616 4333 2621
rect 4340 2616 4345 2621
rect 4351 2616 4356 2621
rect 4363 2616 4368 2621
rect 4374 2616 4379 2621
rect 4394 2606 4398 2612
rect 4404 2606 4408 2612
rect 4419 2589 4423 2615
rect 4429 2589 4433 2615
rect 4444 2595 4448 2615
rect 4454 2595 4458 2615
rect 4464 2595 4468 2615
rect 4474 2595 4478 2615
rect 4484 2595 4488 2615
rect 4494 2595 4498 2615
rect 4504 2605 4508 2615
rect 4519 2515 4523 2615
rect 4529 2515 4533 2615
rect 4539 2515 4543 2615
rect 4549 2515 4553 2615
rect 4559 2515 4563 2615
rect 4569 2515 4573 2615
rect 4579 2560 4583 2615
rect 6311 2637 6316 2642
rect 6322 2637 6327 2642
rect 6349 2637 6354 2642
rect 6360 2637 6365 2642
rect 6376 2637 6381 2642
rect 6387 2637 6392 2642
rect 6399 2637 6404 2642
rect 6410 2637 6415 2642
rect 6422 2637 6427 2642
rect 6433 2637 6438 2642
rect 6453 2627 6457 2633
rect 6463 2627 6467 2633
rect 6478 2610 6482 2636
rect 6488 2610 6492 2636
rect 6503 2616 6507 2636
rect 6513 2616 6517 2636
rect 6523 2616 6527 2636
rect 6533 2616 6537 2636
rect 6543 2616 6547 2636
rect 6553 2616 6557 2636
rect 6563 2626 6567 2636
rect 6578 2536 6582 2636
rect 6588 2536 6592 2636
rect 6598 2536 6602 2636
rect 6608 2536 6612 2636
rect 6618 2536 6622 2636
rect 6628 2536 6632 2636
rect 6638 2581 6642 2636
rect 7989 2775 8092 2791
rect 7989 2492 8092 2508
rect 3349 1911 3452 1927
rect 3349 1628 3452 1644
rect 7989 1929 8092 1945
rect 7989 1646 8092 1662
rect 4597 1055 4601 1110
rect 4607 1055 4611 1155
rect 4617 1055 4621 1155
rect 4627 1055 4631 1155
rect 4637 1055 4641 1155
rect 4647 1055 4651 1155
rect 4657 1055 4661 1155
rect 4672 1055 4676 1065
rect 4682 1055 4686 1075
rect 4692 1055 4696 1075
rect 4702 1055 4706 1075
rect 4712 1055 4716 1075
rect 4722 1055 4726 1075
rect 4732 1055 4736 1075
rect 4747 1055 4751 1081
rect 4757 1055 4761 1081
rect 4772 1058 4776 1064
rect 4782 1058 4786 1064
rect 3349 971 3452 987
rect 3349 688 3452 704
rect 4801 1049 4806 1054
rect 4812 1049 4817 1054
rect 4824 1049 4829 1054
rect 4835 1049 4840 1054
rect 4847 1049 4852 1054
rect 4858 1049 4863 1054
rect 4874 1049 4879 1054
rect 4885 1049 4890 1054
rect 4912 1049 4917 1054
rect 4923 1049 4928 1054
rect 6646 1027 6650 1082
rect 6656 1027 6660 1127
rect 6666 1027 6670 1127
rect 6676 1027 6680 1127
rect 6686 1027 6690 1127
rect 6696 1027 6700 1127
rect 6706 1027 6710 1127
rect 6721 1027 6725 1037
rect 6731 1027 6735 1047
rect 6741 1027 6745 1047
rect 6751 1027 6755 1047
rect 6761 1027 6765 1047
rect 6771 1027 6775 1047
rect 6781 1027 6785 1047
rect 6796 1027 6800 1053
rect 6806 1027 6810 1053
rect 6821 1030 6825 1036
rect 6831 1030 6835 1036
rect 6850 1021 6855 1026
rect 6861 1021 6866 1026
rect 6873 1021 6878 1026
rect 6884 1021 6889 1026
rect 6896 1021 6901 1026
rect 6907 1021 6912 1026
rect 6923 1021 6928 1026
rect 6934 1021 6939 1026
rect 6961 1021 6966 1026
rect 6972 1021 6977 1026
rect 7988 925 8091 941
rect 7988 642 8091 658
rect 3925 -111 3941 -8
rect 4208 -111 4224 -8
rect 5079 -110 5095 -7
rect 5362 -110 5378 -7
rect 6230 -110 6246 -7
rect 6513 -110 6529 -7
rect 7321 -110 7337 -7
rect 7604 -110 7620 -7
<< pdcontact >>
rect 3912 3725 3927 3827
rect 4196 3725 4211 3827
rect 5077 3725 5092 3827
rect 5361 3725 5376 3827
rect 6232 3725 6247 3827
rect 6516 3725 6531 3827
rect 7425 3725 7440 3827
rect 7709 3725 7724 3827
rect 3093 2821 3195 2836
rect 3093 2537 3195 2552
rect 4252 2653 4257 2658
rect 4263 2653 4268 2658
rect 4290 2653 4295 2658
rect 4301 2653 4306 2658
rect 4317 2653 4322 2658
rect 4328 2653 4333 2658
rect 4340 2653 4345 2658
rect 4351 2653 4356 2658
rect 4363 2653 4368 2658
rect 4374 2653 4379 2658
rect 4394 2637 4398 2651
rect 4404 2637 4408 2651
rect 4419 2637 4423 2698
rect 4429 2637 4433 2698
rect 4444 2637 4448 2707
rect 4454 2637 4458 2707
rect 4464 2637 4468 2707
rect 4474 2637 4478 2707
rect 4484 2637 4488 2707
rect 4519 2637 4523 2737
rect 4529 2637 4533 2737
rect 4539 2637 4543 2737
rect 4549 2637 4553 2737
rect 4559 2637 4563 2737
rect 4569 2637 4573 2737
rect 4579 2637 4583 2737
rect 4589 2637 4593 2737
rect 4599 2637 4603 2737
rect 4609 2637 4613 2737
rect 4619 2637 4623 2737
rect 4629 2637 4633 2737
rect 4639 2637 4643 2737
rect 4649 2637 4653 2737
rect 4659 2637 4663 2670
rect 6311 2674 6316 2679
rect 6322 2674 6327 2679
rect 6349 2674 6354 2679
rect 6360 2674 6365 2679
rect 6376 2674 6381 2679
rect 6387 2674 6392 2679
rect 6399 2674 6404 2679
rect 6410 2674 6415 2679
rect 6422 2674 6427 2679
rect 6433 2674 6438 2679
rect 6453 2658 6457 2672
rect 6463 2658 6467 2672
rect 6478 2658 6482 2719
rect 6488 2658 6492 2719
rect 6503 2658 6507 2728
rect 6513 2658 6517 2728
rect 6523 2658 6527 2728
rect 6533 2658 6537 2728
rect 6543 2658 6547 2728
rect 6578 2658 6582 2758
rect 6588 2658 6592 2758
rect 6598 2658 6602 2758
rect 6608 2658 6612 2758
rect 6618 2658 6622 2758
rect 6628 2658 6632 2758
rect 6638 2658 6642 2758
rect 6648 2658 6652 2758
rect 6658 2658 6662 2758
rect 6668 2658 6672 2758
rect 6678 2658 6682 2758
rect 6688 2658 6692 2758
rect 6698 2658 6702 2758
rect 6708 2658 6712 2758
rect 6718 2658 6722 2691
rect 8247 2777 8349 2792
rect 8247 2493 8349 2508
rect 3092 1911 3194 1926
rect 3092 1627 3194 1642
rect 8247 1931 8349 1946
rect 8247 1647 8349 1662
rect 3092 971 3194 986
rect 3092 687 3194 702
rect 4517 1000 4521 1033
rect 4527 933 4531 1033
rect 4537 933 4541 1033
rect 4547 933 4551 1033
rect 4557 933 4561 1033
rect 4567 933 4571 1033
rect 4577 933 4581 1033
rect 4587 933 4591 1033
rect 4597 933 4601 1033
rect 4607 933 4611 1033
rect 4617 933 4621 1033
rect 4627 933 4631 1033
rect 4637 933 4641 1033
rect 4647 933 4651 1033
rect 4657 933 4661 1033
rect 4692 963 4696 1033
rect 4702 963 4706 1033
rect 4712 963 4716 1033
rect 4722 963 4726 1033
rect 4732 963 4736 1033
rect 4747 972 4751 1033
rect 4757 972 4761 1033
rect 4772 1019 4776 1033
rect 4782 1019 4786 1033
rect 4801 1012 4806 1017
rect 4812 1012 4817 1017
rect 4824 1012 4829 1017
rect 4835 1012 4840 1017
rect 4847 1012 4852 1017
rect 4858 1012 4863 1017
rect 4874 1012 4879 1017
rect 4885 1012 4890 1017
rect 4912 1012 4917 1017
rect 4923 1012 4928 1017
rect 6566 972 6570 1005
rect 6576 905 6580 1005
rect 6586 905 6590 1005
rect 6596 905 6600 1005
rect 6606 905 6610 1005
rect 6616 905 6620 1005
rect 6626 905 6630 1005
rect 6636 905 6640 1005
rect 6646 905 6650 1005
rect 6656 905 6660 1005
rect 6666 905 6670 1005
rect 6676 905 6680 1005
rect 6686 905 6690 1005
rect 6696 905 6700 1005
rect 6706 905 6710 1005
rect 6741 935 6745 1005
rect 6751 935 6755 1005
rect 6761 935 6765 1005
rect 6771 935 6775 1005
rect 6781 935 6785 1005
rect 6796 944 6800 1005
rect 6806 944 6810 1005
rect 6821 991 6825 1005
rect 6831 991 6835 1005
rect 6850 984 6855 989
rect 6861 984 6866 989
rect 6873 984 6878 989
rect 6884 984 6889 989
rect 6896 984 6901 989
rect 6907 984 6912 989
rect 6923 984 6928 989
rect 6934 984 6939 989
rect 6961 984 6966 989
rect 6972 984 6977 989
rect 8246 927 8348 942
rect 8246 643 8348 658
rect 3926 -368 3941 -266
rect 4210 -368 4225 -266
rect 5080 -367 5095 -265
rect 5364 -367 5379 -265
rect 6231 -367 6246 -265
rect 6515 -367 6530 -265
rect 7322 -367 7337 -265
rect 7606 -367 7621 -265
<< psubstratepdiff >>
rect 4745 3680 4760 3682
rect 4389 3634 4760 3680
rect 4390 3608 4760 3634
rect 4390 3603 4423 3608
rect 4390 3600 4411 3603
rect 3909 3436 3928 3457
rect 4203 3436 4222 3457
rect 4738 3208 4760 3608
rect 5074 3436 5093 3457
rect 5368 3436 5387 3457
rect 6229 3436 6248 3457
rect 6523 3436 6542 3457
rect 7422 3436 7441 3457
rect 7716 3436 7735 3457
rect 3463 2828 3484 2847
rect 4745 2800 4760 3208
rect 6405 2806 6440 2807
rect 6405 2800 6415 2806
rect 6421 2800 6424 2806
rect 6430 2800 6440 2806
rect 4346 2785 4381 2786
rect 4346 2779 4356 2785
rect 4362 2779 4365 2785
rect 4371 2779 4381 2785
rect 4346 2778 4381 2779
rect 4436 2785 4705 2786
rect 4436 2779 4446 2785
rect 4452 2779 4455 2785
rect 4461 2779 4464 2785
rect 4470 2779 4473 2785
rect 4479 2779 4482 2785
rect 4488 2779 4491 2785
rect 4497 2779 4500 2785
rect 4506 2779 4509 2785
rect 4515 2779 4518 2785
rect 4524 2779 4527 2785
rect 4533 2779 4536 2785
rect 4542 2779 4545 2785
rect 4551 2779 4554 2785
rect 4560 2779 4563 2785
rect 4569 2779 4572 2785
rect 4578 2779 4581 2785
rect 4587 2779 4590 2785
rect 4596 2779 4599 2785
rect 4605 2779 4608 2785
rect 4614 2779 4617 2785
rect 4623 2779 4626 2785
rect 4632 2779 4635 2785
rect 4641 2779 4644 2785
rect 4650 2779 4653 2785
rect 4659 2779 4662 2785
rect 4668 2779 4671 2785
rect 4677 2779 4680 2785
rect 4686 2779 4689 2785
rect 4695 2779 4705 2785
rect 4436 2778 4705 2779
rect 4346 2776 4354 2778
rect 4346 2770 4347 2776
rect 4353 2770 4354 2776
rect 4697 2776 4705 2778
rect 4346 2767 4354 2770
rect 4346 2761 4347 2767
rect 4353 2761 4354 2767
rect 4346 2758 4354 2761
rect 4346 2752 4347 2758
rect 4353 2752 4354 2758
rect 4346 2749 4354 2752
rect 4346 2743 4347 2749
rect 4353 2743 4354 2749
rect 4346 2741 4354 2743
rect 4346 2735 4347 2741
rect 4353 2735 4354 2741
rect 4346 2732 4354 2735
rect 4346 2726 4347 2732
rect 4353 2726 4354 2732
rect 4346 2723 4354 2726
rect 4346 2717 4347 2723
rect 4353 2717 4354 2723
rect 4346 2714 4354 2717
rect 4346 2708 4347 2714
rect 4353 2708 4354 2714
rect 4346 2705 4354 2708
rect 4346 2699 4347 2705
rect 4353 2699 4354 2705
rect 4346 2697 4354 2699
rect 4221 2696 4354 2697
rect 4221 2690 4231 2696
rect 4237 2690 4240 2696
rect 4246 2690 4249 2696
rect 4255 2690 4258 2696
rect 4264 2690 4267 2696
rect 4273 2690 4276 2696
rect 4282 2690 4285 2696
rect 4291 2690 4294 2696
rect 4300 2690 4303 2696
rect 4309 2690 4312 2696
rect 4318 2690 4321 2696
rect 4327 2690 4330 2696
rect 4336 2690 4339 2696
rect 4345 2690 4354 2696
rect 4221 2689 4354 2690
rect 4221 2688 4229 2689
rect 4221 2682 4222 2688
rect 4228 2682 4229 2688
rect 4221 2679 4229 2682
rect 4221 2673 4222 2679
rect 4228 2673 4229 2679
rect 4221 2670 4229 2673
rect 4221 2664 4222 2670
rect 4228 2664 4229 2670
rect 4221 2661 4229 2664
rect 4221 2655 4222 2661
rect 4228 2655 4229 2661
rect 4221 2652 4229 2655
rect 4221 2646 4222 2652
rect 4228 2646 4229 2652
rect 4221 2589 4229 2646
rect 4697 2770 4698 2776
rect 4704 2770 4705 2776
rect 4697 2767 4705 2770
rect 4697 2761 4698 2767
rect 4704 2761 4705 2767
rect 4697 2758 4705 2761
rect 4697 2752 4698 2758
rect 4704 2752 4705 2758
rect 4697 2749 4705 2752
rect 4697 2743 4698 2749
rect 4704 2743 4705 2749
rect 4697 2737 4705 2743
rect 4697 2731 4698 2737
rect 4704 2731 4705 2737
rect 4697 2728 4705 2731
rect 4697 2722 4698 2728
rect 4704 2722 4705 2728
rect 4697 2719 4705 2722
rect 4697 2713 4698 2719
rect 4704 2713 4705 2719
rect 4697 2710 4705 2713
rect 4697 2704 4698 2710
rect 4704 2704 4705 2710
rect 4697 2703 4705 2704
rect 4697 2697 4698 2703
rect 4704 2697 4705 2703
rect 4697 2694 4705 2697
rect 4697 2688 4698 2694
rect 4704 2688 4705 2694
rect 4697 2685 4705 2688
rect 4697 2679 4698 2685
rect 4704 2679 4705 2685
rect 4697 2676 4705 2679
rect 4697 2670 4698 2676
rect 4704 2670 4705 2676
rect 4697 2667 4705 2670
rect 4697 2661 4698 2667
rect 4704 2661 4705 2667
rect 4697 2658 4705 2661
rect 4697 2652 4698 2658
rect 4704 2652 4705 2658
rect 4697 2615 4705 2652
rect 4745 2631 4757 2800
rect 6405 2799 6440 2800
rect 6495 2806 6764 2807
rect 6495 2800 6505 2806
rect 6511 2800 6514 2806
rect 6520 2800 6523 2806
rect 6529 2800 6532 2806
rect 6538 2800 6541 2806
rect 6547 2800 6550 2806
rect 6556 2800 6559 2806
rect 6565 2800 6568 2806
rect 6574 2800 6577 2806
rect 6583 2800 6586 2806
rect 6592 2800 6595 2806
rect 6601 2800 6604 2806
rect 6610 2800 6613 2806
rect 6619 2800 6622 2806
rect 6628 2800 6631 2806
rect 6637 2800 6640 2806
rect 6646 2800 6649 2806
rect 6655 2800 6658 2806
rect 6664 2800 6667 2806
rect 6673 2800 6676 2806
rect 6682 2800 6685 2806
rect 6691 2800 6694 2806
rect 6700 2800 6703 2806
rect 6709 2800 6712 2806
rect 6718 2800 6721 2806
rect 6727 2800 6730 2806
rect 6736 2800 6739 2806
rect 6745 2800 6748 2806
rect 6754 2800 6764 2806
rect 6495 2799 6764 2800
rect 6405 2797 6413 2799
rect 6405 2791 6406 2797
rect 6412 2791 6413 2797
rect 6756 2797 6764 2799
rect 6405 2788 6413 2791
rect 6405 2782 6406 2788
rect 6412 2782 6413 2788
rect 6405 2779 6413 2782
rect 6405 2773 6406 2779
rect 6412 2773 6413 2779
rect 6405 2770 6413 2773
rect 6405 2764 6406 2770
rect 6412 2764 6413 2770
rect 6405 2762 6413 2764
rect 6405 2756 6406 2762
rect 6412 2756 6413 2762
rect 6405 2753 6413 2756
rect 6405 2747 6406 2753
rect 6412 2747 6413 2753
rect 6405 2744 6413 2747
rect 6405 2738 6406 2744
rect 6412 2738 6413 2744
rect 6405 2735 6413 2738
rect 6405 2729 6406 2735
rect 6412 2729 6413 2735
rect 6405 2726 6413 2729
rect 6405 2720 6406 2726
rect 6412 2720 6413 2726
rect 6405 2718 6413 2720
rect 4708 2626 4757 2631
rect 6280 2717 6413 2718
rect 6280 2711 6290 2717
rect 6296 2711 6299 2717
rect 6305 2711 6308 2717
rect 6314 2711 6317 2717
rect 6323 2711 6326 2717
rect 6332 2711 6335 2717
rect 6341 2711 6344 2717
rect 6350 2711 6353 2717
rect 6359 2711 6362 2717
rect 6368 2711 6371 2717
rect 6377 2711 6380 2717
rect 6386 2711 6389 2717
rect 6395 2711 6398 2717
rect 6404 2711 6413 2717
rect 6280 2710 6413 2711
rect 6280 2709 6288 2710
rect 6280 2703 6281 2709
rect 6287 2703 6288 2709
rect 6280 2700 6288 2703
rect 6280 2694 6281 2700
rect 6287 2694 6288 2700
rect 6280 2691 6288 2694
rect 6280 2685 6281 2691
rect 6287 2685 6288 2691
rect 6280 2682 6288 2685
rect 6280 2676 6281 2682
rect 6287 2676 6288 2682
rect 6280 2673 6288 2676
rect 6280 2667 6281 2673
rect 6287 2667 6288 2673
rect 4221 2583 4222 2589
rect 4228 2583 4229 2589
rect 4221 2582 4229 2583
rect 4221 2581 4369 2582
rect 4221 2575 4231 2581
rect 4237 2575 4240 2581
rect 4246 2575 4249 2581
rect 4255 2575 4258 2581
rect 4264 2575 4267 2581
rect 4273 2575 4276 2581
rect 4282 2575 4285 2581
rect 4291 2575 4294 2581
rect 4300 2575 4303 2581
rect 4309 2575 4312 2581
rect 4318 2575 4321 2581
rect 4327 2575 4330 2581
rect 4336 2575 4339 2581
rect 4345 2575 4348 2581
rect 4354 2575 4355 2581
rect 4361 2575 4369 2581
rect 4221 2574 4369 2575
rect 3463 2534 3484 2553
rect 4361 2572 4369 2574
rect 4361 2566 4362 2572
rect 4368 2566 4369 2572
rect 4361 2563 4369 2566
rect 4361 2557 4362 2563
rect 4368 2557 4369 2563
rect 4361 2556 4475 2557
rect 4361 2550 4371 2556
rect 4377 2550 4380 2556
rect 4386 2550 4389 2556
rect 4395 2550 4398 2556
rect 4404 2550 4407 2556
rect 4413 2550 4416 2556
rect 4422 2550 4425 2556
rect 4431 2550 4434 2556
rect 4440 2550 4443 2556
rect 4449 2550 4452 2556
rect 4458 2550 4461 2556
rect 4467 2550 4475 2556
rect 4361 2549 4475 2550
rect 4467 2547 4475 2549
rect 4467 2541 4468 2547
rect 4474 2541 4475 2547
rect 4467 2538 4475 2541
rect 4467 2532 4468 2538
rect 4474 2532 4475 2538
rect 4467 2529 4475 2532
rect 4467 2523 4468 2529
rect 4474 2523 4475 2529
rect 4467 2520 4475 2523
rect 4467 2514 4468 2520
rect 4474 2514 4475 2520
rect 4599 2614 4705 2615
rect 4599 2608 4609 2614
rect 4615 2608 4618 2614
rect 4624 2608 4627 2614
rect 4633 2608 4636 2614
rect 4642 2608 4645 2614
rect 4651 2608 4654 2614
rect 4660 2608 4663 2614
rect 4669 2608 4672 2614
rect 4678 2608 4681 2614
rect 4687 2608 4690 2614
rect 4696 2608 4705 2614
rect 4599 2607 4705 2608
rect 6280 2610 6288 2667
rect 6756 2791 6757 2797
rect 6763 2791 6764 2797
rect 6756 2788 6764 2791
rect 6756 2782 6757 2788
rect 6763 2782 6764 2788
rect 6756 2779 6764 2782
rect 6756 2773 6757 2779
rect 6763 2773 6764 2779
rect 6756 2770 6764 2773
rect 6756 2764 6757 2770
rect 6763 2764 6764 2770
rect 6756 2758 6764 2764
rect 6756 2752 6757 2758
rect 6763 2752 6764 2758
rect 6756 2749 6764 2752
rect 6756 2743 6757 2749
rect 6763 2743 6764 2749
rect 6756 2740 6764 2743
rect 6756 2734 6757 2740
rect 6763 2734 6764 2740
rect 6756 2731 6764 2734
rect 6756 2725 6757 2731
rect 6763 2725 6764 2731
rect 6756 2724 6764 2725
rect 6756 2718 6757 2724
rect 6763 2718 6764 2724
rect 6756 2715 6764 2718
rect 6756 2709 6757 2715
rect 6763 2709 6764 2715
rect 6756 2706 6764 2709
rect 6756 2700 6757 2706
rect 6763 2700 6764 2706
rect 6756 2697 6764 2700
rect 6756 2691 6757 2697
rect 6763 2691 6764 2697
rect 6756 2688 6764 2691
rect 6756 2682 6757 2688
rect 6763 2682 6764 2688
rect 6756 2679 6764 2682
rect 6756 2673 6757 2679
rect 6763 2673 6764 2679
rect 6756 2636 6764 2673
rect 4599 2605 4607 2607
rect 4599 2599 4600 2605
rect 4606 2599 4607 2605
rect 4599 2596 4607 2599
rect 4599 2590 4600 2596
rect 4606 2590 4607 2596
rect 6280 2604 6281 2610
rect 6287 2604 6288 2610
rect 6280 2603 6288 2604
rect 6280 2602 6428 2603
rect 6280 2596 6290 2602
rect 6296 2596 6299 2602
rect 6305 2596 6308 2602
rect 6314 2596 6317 2602
rect 6323 2596 6326 2602
rect 6332 2596 6335 2602
rect 6341 2596 6344 2602
rect 6350 2596 6353 2602
rect 6359 2596 6362 2602
rect 6368 2596 6371 2602
rect 6377 2596 6380 2602
rect 6386 2596 6389 2602
rect 6395 2596 6398 2602
rect 6404 2596 6407 2602
rect 6413 2596 6414 2602
rect 6420 2596 6428 2602
rect 6280 2595 6428 2596
rect 4599 2587 4607 2590
rect 4599 2581 4600 2587
rect 4606 2581 4607 2587
rect 4599 2578 4607 2581
rect 4599 2572 4600 2578
rect 4606 2572 4607 2578
rect 4599 2569 4607 2572
rect 6420 2593 6428 2595
rect 6420 2587 6421 2593
rect 6427 2587 6428 2593
rect 6420 2584 6428 2587
rect 6420 2578 6421 2584
rect 6427 2578 6428 2584
rect 6420 2577 6534 2578
rect 6420 2571 6430 2577
rect 6436 2571 6439 2577
rect 6445 2571 6448 2577
rect 6454 2571 6457 2577
rect 6463 2571 6466 2577
rect 6472 2571 6475 2577
rect 6481 2571 6484 2577
rect 6490 2571 6493 2577
rect 6499 2571 6502 2577
rect 6508 2571 6511 2577
rect 6517 2571 6520 2577
rect 6526 2571 6534 2577
rect 6420 2570 6534 2571
rect 4599 2563 4600 2569
rect 4606 2563 4607 2569
rect 4599 2560 4607 2563
rect 4599 2554 4600 2560
rect 4606 2554 4607 2560
rect 4599 2551 4607 2554
rect 4599 2545 4600 2551
rect 4606 2545 4607 2551
rect 4599 2542 4607 2545
rect 4599 2536 4600 2542
rect 4606 2536 4607 2542
rect 4599 2533 4607 2536
rect 4599 2527 4600 2533
rect 4606 2527 4607 2533
rect 4599 2524 4607 2527
rect 4599 2518 4600 2524
rect 4606 2518 4607 2524
rect 4599 2515 4607 2518
rect 4467 2511 4475 2514
rect 4467 2505 4468 2511
rect 4474 2505 4475 2511
rect 4467 2502 4475 2505
rect 4467 2496 4468 2502
rect 4474 2496 4475 2502
rect 4467 2491 4475 2496
rect 4599 2509 4600 2515
rect 4606 2509 4607 2515
rect 4599 2506 4607 2509
rect 4599 2500 4600 2506
rect 4606 2500 4607 2506
rect 6526 2568 6534 2570
rect 6526 2562 6527 2568
rect 6533 2562 6534 2568
rect 6526 2559 6534 2562
rect 6526 2553 6527 2559
rect 6533 2553 6534 2559
rect 6526 2550 6534 2553
rect 6526 2544 6527 2550
rect 6533 2544 6534 2550
rect 6526 2541 6534 2544
rect 6526 2535 6527 2541
rect 6533 2535 6534 2541
rect 6658 2635 6764 2636
rect 6658 2629 6668 2635
rect 6674 2629 6677 2635
rect 6683 2629 6686 2635
rect 6692 2629 6695 2635
rect 6701 2629 6704 2635
rect 6710 2629 6713 2635
rect 6719 2629 6722 2635
rect 6728 2629 6731 2635
rect 6737 2629 6740 2635
rect 6746 2629 6749 2635
rect 6755 2629 6764 2635
rect 6658 2628 6764 2629
rect 7958 2776 7979 2795
rect 6658 2626 6666 2628
rect 6658 2620 6659 2626
rect 6665 2620 6666 2626
rect 6658 2617 6666 2620
rect 6658 2611 6659 2617
rect 6665 2611 6666 2617
rect 6658 2608 6666 2611
rect 6658 2602 6659 2608
rect 6665 2602 6666 2608
rect 6658 2599 6666 2602
rect 6658 2593 6659 2599
rect 6665 2593 6666 2599
rect 6658 2590 6666 2593
rect 6658 2584 6659 2590
rect 6665 2584 6666 2590
rect 6658 2581 6666 2584
rect 6658 2575 6659 2581
rect 6665 2575 6666 2581
rect 6658 2572 6666 2575
rect 6658 2566 6659 2572
rect 6665 2566 6666 2572
rect 6658 2563 6666 2566
rect 6658 2557 6659 2563
rect 6665 2557 6666 2563
rect 6658 2554 6666 2557
rect 6658 2548 6659 2554
rect 6665 2548 6666 2554
rect 6658 2545 6666 2548
rect 6658 2539 6659 2545
rect 6665 2539 6666 2545
rect 6658 2536 6666 2539
rect 6526 2532 6534 2535
rect 6526 2526 6527 2532
rect 6533 2526 6534 2532
rect 6526 2523 6534 2526
rect 6526 2517 6527 2523
rect 6533 2517 6534 2523
rect 6526 2512 6534 2517
rect 6658 2530 6659 2536
rect 6665 2530 6666 2536
rect 6658 2527 6666 2530
rect 6658 2521 6659 2527
rect 6665 2521 6666 2527
rect 6658 2518 6666 2521
rect 6658 2512 6659 2518
rect 6665 2512 6666 2518
rect 6526 2511 6666 2512
rect 6526 2505 6536 2511
rect 6542 2505 6545 2511
rect 6551 2505 6554 2511
rect 6560 2505 6563 2511
rect 6569 2505 6572 2511
rect 6578 2505 6581 2511
rect 6587 2505 6590 2511
rect 6596 2505 6599 2511
rect 6605 2505 6608 2511
rect 6614 2505 6617 2511
rect 6623 2505 6626 2511
rect 6632 2505 6635 2511
rect 6641 2505 6644 2511
rect 6650 2505 6653 2511
rect 6659 2505 6666 2511
rect 6526 2504 6666 2505
rect 4599 2497 4607 2500
rect 4599 2491 4600 2497
rect 4606 2491 4607 2497
rect 4467 2490 4607 2491
rect 4467 2484 4477 2490
rect 4483 2484 4486 2490
rect 4492 2484 4495 2490
rect 4501 2484 4504 2490
rect 4510 2484 4513 2490
rect 4519 2484 4522 2490
rect 4528 2484 4531 2490
rect 4537 2484 4540 2490
rect 4546 2484 4549 2490
rect 4555 2484 4558 2490
rect 4564 2484 4567 2490
rect 4573 2484 4576 2490
rect 4582 2484 4585 2490
rect 4591 2484 4594 2490
rect 4600 2484 4607 2490
rect 4467 2483 4607 2484
rect 7958 2482 7979 2501
rect 3462 1918 3483 1937
rect 3462 1624 3483 1643
rect 7958 1930 7979 1949
rect 7958 1636 7979 1655
rect 4573 1186 4713 1187
rect 4573 1180 4580 1186
rect 4586 1180 4589 1186
rect 4595 1180 4598 1186
rect 4604 1180 4607 1186
rect 4613 1180 4616 1186
rect 4622 1180 4625 1186
rect 4631 1180 4634 1186
rect 4640 1180 4643 1186
rect 4649 1180 4652 1186
rect 4658 1180 4661 1186
rect 4667 1180 4670 1186
rect 4676 1180 4679 1186
rect 4685 1180 4688 1186
rect 4694 1180 4697 1186
rect 4703 1180 4713 1186
rect 4573 1179 4713 1180
rect 4573 1173 4574 1179
rect 4580 1173 4581 1179
rect 4573 1170 4581 1173
rect 4573 1164 4574 1170
rect 4580 1164 4581 1170
rect 4573 1161 4581 1164
rect 4573 1155 4574 1161
rect 4580 1155 4581 1161
rect 4705 1174 4713 1179
rect 4705 1168 4706 1174
rect 4712 1168 4713 1174
rect 4705 1165 4713 1168
rect 4705 1159 4706 1165
rect 4712 1159 4713 1165
rect 4705 1156 4713 1159
rect 4573 1152 4581 1155
rect 4573 1146 4574 1152
rect 4580 1146 4581 1152
rect 4573 1143 4581 1146
rect 4573 1137 4574 1143
rect 4580 1137 4581 1143
rect 4573 1134 4581 1137
rect 4573 1128 4574 1134
rect 4580 1128 4581 1134
rect 4573 1125 4581 1128
rect 4573 1119 4574 1125
rect 4580 1119 4581 1125
rect 4573 1116 4581 1119
rect 4573 1110 4574 1116
rect 4580 1110 4581 1116
rect 4573 1107 4581 1110
rect 4573 1101 4574 1107
rect 4580 1101 4581 1107
rect 4573 1098 4581 1101
rect 4573 1092 4574 1098
rect 4580 1092 4581 1098
rect 4573 1089 4581 1092
rect 4573 1083 4574 1089
rect 4580 1083 4581 1089
rect 4573 1080 4581 1083
rect 4573 1074 4574 1080
rect 4580 1074 4581 1080
rect 4573 1071 4581 1074
rect 4573 1065 4574 1071
rect 4580 1065 4581 1071
rect 4573 1063 4581 1065
rect 4475 1062 4581 1063
rect 4475 1056 4484 1062
rect 4490 1056 4493 1062
rect 4499 1056 4502 1062
rect 4508 1056 4511 1062
rect 4517 1056 4520 1062
rect 4526 1056 4529 1062
rect 4535 1056 4538 1062
rect 4544 1056 4547 1062
rect 4553 1056 4556 1062
rect 4562 1056 4565 1062
rect 4571 1056 4581 1062
rect 4475 1055 4581 1056
rect 4705 1150 4706 1156
rect 4712 1150 4713 1156
rect 4705 1147 4713 1150
rect 4705 1141 4706 1147
rect 4712 1141 4713 1147
rect 4705 1138 4713 1141
rect 4705 1132 4706 1138
rect 4712 1132 4713 1138
rect 4705 1129 4713 1132
rect 4705 1123 4706 1129
rect 4712 1123 4713 1129
rect 4705 1121 4713 1123
rect 6622 1158 6762 1159
rect 6622 1152 6629 1158
rect 6635 1152 6638 1158
rect 6644 1152 6647 1158
rect 6653 1152 6656 1158
rect 6662 1152 6665 1158
rect 6671 1152 6674 1158
rect 6680 1152 6683 1158
rect 6689 1152 6692 1158
rect 6698 1152 6701 1158
rect 6707 1152 6710 1158
rect 6716 1152 6719 1158
rect 6725 1152 6728 1158
rect 6734 1152 6737 1158
rect 6743 1152 6746 1158
rect 6752 1152 6762 1158
rect 6622 1151 6762 1152
rect 6622 1145 6623 1151
rect 6629 1145 6630 1151
rect 6622 1142 6630 1145
rect 6622 1136 6623 1142
rect 6629 1136 6630 1142
rect 6622 1133 6630 1136
rect 6622 1127 6623 1133
rect 6629 1127 6630 1133
rect 6754 1146 6762 1151
rect 6754 1140 6755 1146
rect 6761 1140 6762 1146
rect 6754 1137 6762 1140
rect 6754 1131 6755 1137
rect 6761 1131 6762 1137
rect 6754 1128 6762 1131
rect 6622 1124 6630 1127
rect 4705 1120 4819 1121
rect 4705 1114 4713 1120
rect 4719 1114 4722 1120
rect 4728 1114 4731 1120
rect 4737 1114 4740 1120
rect 4746 1114 4749 1120
rect 4755 1114 4758 1120
rect 4764 1114 4767 1120
rect 4773 1114 4776 1120
rect 4782 1114 4785 1120
rect 4791 1114 4794 1120
rect 4800 1114 4803 1120
rect 4809 1114 4819 1120
rect 4705 1113 4819 1114
rect 4811 1107 4812 1113
rect 4818 1107 4819 1113
rect 4811 1104 4819 1107
rect 4811 1098 4812 1104
rect 4818 1098 4819 1104
rect 4811 1096 4819 1098
rect 6622 1118 6623 1124
rect 6629 1118 6630 1124
rect 6622 1115 6630 1118
rect 6622 1109 6623 1115
rect 6629 1109 6630 1115
rect 6622 1106 6630 1109
rect 6622 1100 6623 1106
rect 6629 1100 6630 1106
rect 6622 1097 6630 1100
rect 4811 1095 4959 1096
rect 4811 1089 4819 1095
rect 4825 1089 4826 1095
rect 4832 1089 4835 1095
rect 4841 1089 4844 1095
rect 4850 1089 4853 1095
rect 4859 1089 4862 1095
rect 4868 1089 4871 1095
rect 4877 1089 4880 1095
rect 4886 1089 4889 1095
rect 4895 1089 4898 1095
rect 4904 1089 4907 1095
rect 4913 1089 4916 1095
rect 4922 1089 4925 1095
rect 4931 1089 4934 1095
rect 4940 1089 4943 1095
rect 4949 1089 4959 1095
rect 4811 1088 4959 1089
rect 4951 1087 4959 1088
rect 4951 1081 4952 1087
rect 4958 1081 4959 1087
rect 3462 978 3483 997
rect 4475 1018 4483 1055
rect 4475 1012 4476 1018
rect 4482 1012 4483 1018
rect 4475 1009 4483 1012
rect 4475 1003 4476 1009
rect 4482 1003 4483 1009
rect 4475 1000 4483 1003
rect 4475 994 4476 1000
rect 4482 994 4483 1000
rect 4475 991 4483 994
rect 4475 985 4476 991
rect 4482 985 4483 991
rect 4475 982 4483 985
rect 4475 976 4476 982
rect 4482 976 4483 982
rect 4475 973 4483 976
rect 4475 967 4476 973
rect 4482 967 4483 973
rect 4475 966 4483 967
rect 4475 960 4476 966
rect 4482 960 4483 966
rect 4475 957 4483 960
rect 4475 951 4476 957
rect 4482 951 4483 957
rect 4475 948 4483 951
rect 4475 942 4476 948
rect 4482 942 4483 948
rect 4475 939 4483 942
rect 4475 933 4476 939
rect 4482 933 4483 939
rect 4475 927 4483 933
rect 4475 921 4476 927
rect 4482 921 4483 927
rect 4475 918 4483 921
rect 4475 912 4476 918
rect 4482 912 4483 918
rect 4475 909 4483 912
rect 4475 903 4476 909
rect 4482 903 4483 909
rect 4475 900 4483 903
rect 4475 894 4476 900
rect 4482 894 4483 900
rect 4951 1024 4959 1081
rect 6622 1091 6623 1097
rect 6629 1091 6630 1097
rect 6622 1088 6630 1091
rect 6622 1082 6623 1088
rect 6629 1082 6630 1088
rect 6622 1079 6630 1082
rect 6622 1073 6623 1079
rect 6629 1073 6630 1079
rect 6622 1070 6630 1073
rect 6622 1064 6623 1070
rect 6629 1064 6630 1070
rect 6622 1061 6630 1064
rect 6622 1055 6623 1061
rect 6629 1055 6630 1061
rect 6622 1052 6630 1055
rect 6622 1046 6623 1052
rect 6629 1046 6630 1052
rect 6622 1043 6630 1046
rect 6622 1037 6623 1043
rect 6629 1037 6630 1043
rect 6622 1035 6630 1037
rect 4951 1018 4952 1024
rect 4958 1018 4959 1024
rect 4951 1015 4959 1018
rect 4951 1009 4952 1015
rect 4958 1009 4959 1015
rect 4951 1006 4959 1009
rect 4951 1000 4952 1006
rect 4958 1000 4959 1006
rect 4951 997 4959 1000
rect 4951 991 4952 997
rect 4958 991 4959 997
rect 4951 988 4959 991
rect 4951 982 4952 988
rect 4958 982 4959 988
rect 4951 981 4959 982
rect 4826 980 4959 981
rect 4826 974 4835 980
rect 4841 974 4844 980
rect 4850 974 4853 980
rect 4859 974 4862 980
rect 4868 974 4871 980
rect 4877 974 4880 980
rect 4886 974 4889 980
rect 4895 974 4898 980
rect 4904 974 4907 980
rect 4913 974 4916 980
rect 4922 974 4925 980
rect 4931 974 4934 980
rect 4940 974 4943 980
rect 4949 974 4959 980
rect 4826 973 4959 974
rect 6524 1034 6630 1035
rect 6524 1028 6533 1034
rect 6539 1028 6542 1034
rect 6548 1028 6551 1034
rect 6557 1028 6560 1034
rect 6566 1028 6569 1034
rect 6575 1028 6578 1034
rect 6584 1028 6587 1034
rect 6593 1028 6596 1034
rect 6602 1028 6605 1034
rect 6611 1028 6614 1034
rect 6620 1028 6630 1034
rect 6524 1027 6630 1028
rect 6754 1122 6755 1128
rect 6761 1122 6762 1128
rect 6754 1119 6762 1122
rect 6754 1113 6755 1119
rect 6761 1113 6762 1119
rect 6754 1110 6762 1113
rect 6754 1104 6755 1110
rect 6761 1104 6762 1110
rect 6754 1101 6762 1104
rect 6754 1095 6755 1101
rect 6761 1095 6762 1101
rect 6754 1093 6762 1095
rect 6754 1092 6868 1093
rect 6754 1086 6762 1092
rect 6768 1086 6771 1092
rect 6777 1086 6780 1092
rect 6786 1086 6789 1092
rect 6795 1086 6798 1092
rect 6804 1086 6807 1092
rect 6813 1086 6816 1092
rect 6822 1086 6825 1092
rect 6831 1086 6834 1092
rect 6840 1086 6843 1092
rect 6849 1086 6852 1092
rect 6858 1086 6868 1092
rect 6754 1085 6868 1086
rect 6860 1079 6861 1085
rect 6867 1079 6868 1085
rect 6860 1076 6868 1079
rect 6860 1070 6861 1076
rect 6867 1070 6868 1076
rect 6860 1068 6868 1070
rect 6860 1067 7008 1068
rect 6860 1061 6868 1067
rect 6874 1061 6875 1067
rect 6881 1061 6884 1067
rect 6890 1061 6893 1067
rect 6899 1061 6902 1067
rect 6908 1061 6911 1067
rect 6917 1061 6920 1067
rect 6926 1061 6929 1067
rect 6935 1061 6938 1067
rect 6944 1061 6947 1067
rect 6953 1061 6956 1067
rect 6962 1061 6965 1067
rect 6971 1061 6974 1067
rect 6980 1061 6983 1067
rect 6989 1061 6992 1067
rect 6998 1061 7008 1067
rect 6860 1060 7008 1061
rect 7000 1059 7008 1060
rect 7000 1053 7001 1059
rect 7007 1053 7008 1059
rect 6524 990 6532 1027
rect 6524 984 6525 990
rect 6531 984 6532 990
rect 6524 981 6532 984
rect 6524 975 6525 981
rect 6531 975 6532 981
rect 4826 971 4834 973
rect 4826 965 4827 971
rect 4833 965 4834 971
rect 4826 962 4834 965
rect 4826 956 4827 962
rect 4833 956 4834 962
rect 4826 953 4834 956
rect 4826 947 4827 953
rect 4833 947 4834 953
rect 4826 944 4834 947
rect 4826 938 4827 944
rect 4833 938 4834 944
rect 4826 935 4834 938
rect 4826 929 4827 935
rect 4833 929 4834 935
rect 4826 927 4834 929
rect 4826 921 4827 927
rect 4833 921 4834 927
rect 4826 918 4834 921
rect 4826 912 4827 918
rect 4833 912 4834 918
rect 4826 909 4834 912
rect 4826 903 4827 909
rect 4833 903 4834 909
rect 4826 900 4834 903
rect 4475 892 4483 894
rect 4826 894 4827 900
rect 4833 894 4834 900
rect 4826 892 4834 894
rect 4475 891 4744 892
rect 4475 885 4485 891
rect 4491 885 4494 891
rect 4500 885 4503 891
rect 4509 885 4512 891
rect 4518 885 4521 891
rect 4527 885 4530 891
rect 4536 885 4539 891
rect 4545 885 4548 891
rect 4554 885 4557 891
rect 4563 885 4566 891
rect 4572 885 4575 891
rect 4581 885 4584 891
rect 4590 885 4593 891
rect 4599 885 4602 891
rect 4608 885 4611 891
rect 4617 885 4620 891
rect 4626 885 4629 891
rect 4635 885 4638 891
rect 4644 885 4647 891
rect 4653 885 4656 891
rect 4662 885 4665 891
rect 4671 885 4674 891
rect 4680 885 4683 891
rect 4689 885 4692 891
rect 4698 885 4701 891
rect 4707 885 4710 891
rect 4716 885 4719 891
rect 4725 885 4728 891
rect 4734 885 4744 891
rect 4475 884 4744 885
rect 4799 891 4834 892
rect 4799 885 4809 891
rect 4815 885 4818 891
rect 4824 885 4834 891
rect 4799 884 4834 885
rect 6524 972 6532 975
rect 6524 966 6525 972
rect 6531 966 6532 972
rect 6524 963 6532 966
rect 6524 957 6525 963
rect 6531 957 6532 963
rect 6524 954 6532 957
rect 6524 948 6525 954
rect 6531 948 6532 954
rect 6524 945 6532 948
rect 6524 939 6525 945
rect 6531 939 6532 945
rect 6524 938 6532 939
rect 6524 932 6525 938
rect 6531 932 6532 938
rect 6524 929 6532 932
rect 6524 923 6525 929
rect 6531 923 6532 929
rect 6524 920 6532 923
rect 6524 914 6525 920
rect 6531 914 6532 920
rect 6524 911 6532 914
rect 6524 905 6525 911
rect 6531 905 6532 911
rect 6524 899 6532 905
rect 6524 893 6525 899
rect 6531 893 6532 899
rect 6524 890 6532 893
rect 6524 884 6525 890
rect 6531 884 6532 890
rect 6524 881 6532 884
rect 6524 875 6525 881
rect 6531 875 6532 881
rect 6524 872 6532 875
rect 6524 866 6525 872
rect 6531 866 6532 872
rect 7000 996 7008 1053
rect 7831 1043 7866 1266
rect 7081 1042 7866 1043
rect 7078 1041 7866 1042
rect 7075 1039 7866 1041
rect 7020 1038 7866 1039
rect 7017 1032 7866 1038
rect 7592 1008 7866 1019
rect 7000 990 7001 996
rect 7007 990 7008 996
rect 7000 987 7008 990
rect 7000 981 7001 987
rect 7007 981 7008 987
rect 7000 978 7008 981
rect 7000 972 7001 978
rect 7007 972 7008 978
rect 7000 969 7008 972
rect 7000 963 7001 969
rect 7007 963 7008 969
rect 7000 960 7008 963
rect 7000 954 7001 960
rect 7007 954 7008 960
rect 7000 953 7008 954
rect 6875 952 7008 953
rect 6875 946 6884 952
rect 6890 946 6893 952
rect 6899 946 6902 952
rect 6908 946 6911 952
rect 6917 946 6920 952
rect 6926 946 6929 952
rect 6935 946 6938 952
rect 6944 946 6947 952
rect 6953 946 6956 952
rect 6962 946 6965 952
rect 6971 946 6974 952
rect 6980 946 6983 952
rect 6989 946 6992 952
rect 6998 946 7008 952
rect 6875 945 7008 946
rect 6875 943 6883 945
rect 6875 937 6876 943
rect 6882 937 6883 943
rect 6875 934 6883 937
rect 6875 928 6876 934
rect 6882 928 6883 934
rect 6875 925 6883 928
rect 6875 919 6876 925
rect 6882 919 6883 925
rect 6875 916 6883 919
rect 6875 910 6876 916
rect 6882 910 6883 916
rect 6875 907 6883 910
rect 6875 901 6876 907
rect 6882 901 6883 907
rect 6875 899 6883 901
rect 6875 893 6876 899
rect 6882 893 6883 899
rect 6875 890 6883 893
rect 6875 884 6876 890
rect 6882 884 6883 890
rect 6875 881 6883 884
rect 6875 875 6876 881
rect 6882 875 6883 881
rect 6875 872 6883 875
rect 6524 864 6532 866
rect 6875 866 6876 872
rect 6882 866 6883 872
rect 6875 864 6883 866
rect 6524 863 6793 864
rect 6524 857 6534 863
rect 6540 857 6543 863
rect 6549 857 6552 863
rect 6558 857 6561 863
rect 6567 857 6570 863
rect 6576 857 6579 863
rect 6585 857 6588 863
rect 6594 857 6597 863
rect 6603 857 6606 863
rect 6612 857 6615 863
rect 6621 857 6624 863
rect 6630 857 6633 863
rect 6639 857 6642 863
rect 6648 857 6651 863
rect 6657 857 6660 863
rect 6666 857 6669 863
rect 6675 857 6678 863
rect 6684 857 6687 863
rect 6693 857 6696 863
rect 6702 857 6705 863
rect 6711 857 6714 863
rect 6720 857 6723 863
rect 6729 857 6732 863
rect 6738 857 6741 863
rect 6747 857 6750 863
rect 6756 857 6759 863
rect 6765 857 6768 863
rect 6774 857 6777 863
rect 6783 857 6793 863
rect 6524 856 6793 857
rect 6848 863 6883 864
rect 6848 857 6849 863
rect 6855 857 6858 863
rect 6864 857 6867 863
rect 6873 857 6883 863
rect 6848 856 6883 857
rect 7957 926 7978 945
rect 3462 684 3483 703
rect 7957 632 7978 651
rect 3915 2 3934 23
rect 4209 2 4228 23
rect 5069 3 5088 24
rect 5363 3 5382 24
rect 6220 3 6239 24
rect 6514 3 6533 24
rect 7311 3 7330 24
rect 7605 3 7624 24
<< nsubstratendiff >>
rect 3907 3831 3930 3850
rect 4195 3831 4220 3850
rect 5072 3831 5095 3850
rect 5360 3831 5385 3850
rect 6227 3831 6250 3850
rect 6515 3831 6540 3850
rect 7420 3831 7443 3850
rect 7708 3831 7733 3850
rect 3070 2820 3089 2845
rect 3070 2532 3089 2555
rect 4365 2771 4687 2772
rect 4365 2765 4375 2771
rect 4381 2765 4384 2771
rect 4390 2765 4393 2771
rect 4399 2765 4402 2771
rect 4408 2765 4413 2771
rect 4419 2765 4422 2771
rect 4428 2765 4431 2771
rect 4437 2765 4440 2771
rect 4446 2765 4449 2771
rect 4455 2765 4460 2771
rect 4466 2765 4469 2771
rect 4475 2765 4478 2771
rect 4484 2765 4487 2771
rect 4493 2765 4496 2771
rect 4502 2765 4505 2771
rect 4511 2765 4514 2771
rect 4520 2765 4523 2771
rect 4529 2765 4532 2771
rect 4538 2765 4543 2771
rect 4549 2765 4552 2771
rect 4558 2765 4561 2771
rect 4567 2765 4570 2771
rect 4576 2765 4579 2771
rect 4585 2765 4590 2771
rect 4596 2765 4599 2771
rect 4605 2765 4608 2771
rect 4614 2765 4617 2771
rect 4623 2765 4626 2771
rect 4632 2765 4635 2771
rect 4641 2765 4644 2771
rect 4650 2765 4653 2771
rect 4659 2765 4662 2771
rect 4668 2765 4671 2771
rect 4677 2765 4687 2771
rect 4365 2764 4687 2765
rect 4365 2762 4373 2764
rect 4365 2756 4366 2762
rect 4372 2756 4373 2762
rect 4365 2753 4373 2756
rect 4365 2747 4366 2753
rect 4372 2747 4373 2753
rect 4365 2744 4373 2747
rect 4365 2738 4366 2744
rect 4372 2738 4373 2744
rect 4679 2762 4687 2764
rect 4679 2756 4680 2762
rect 4686 2756 4687 2762
rect 4679 2753 4687 2756
rect 4679 2747 4680 2753
rect 4686 2747 4687 2753
rect 4679 2744 4687 2747
rect 4365 2735 4373 2738
rect 4679 2738 4680 2744
rect 4686 2738 4687 2744
rect 4365 2729 4366 2735
rect 4372 2729 4373 2735
rect 4365 2727 4373 2729
rect 4365 2721 4366 2727
rect 4372 2721 4373 2727
rect 4365 2718 4373 2721
rect 4365 2712 4366 2718
rect 4372 2712 4373 2718
rect 4365 2709 4373 2712
rect 4365 2703 4366 2709
rect 4372 2703 4373 2709
rect 4365 2700 4373 2703
rect 4365 2694 4366 2700
rect 4372 2694 4373 2700
rect 4365 2691 4373 2694
rect 4365 2685 4366 2691
rect 4372 2685 4373 2691
rect 4365 2683 4373 2685
rect 4235 2682 4373 2683
rect 4235 2676 4245 2682
rect 4251 2676 4254 2682
rect 4260 2676 4263 2682
rect 4269 2676 4272 2682
rect 4278 2676 4283 2682
rect 4289 2676 4292 2682
rect 4298 2676 4301 2682
rect 4307 2676 4310 2682
rect 4316 2676 4319 2682
rect 4325 2676 4330 2682
rect 4336 2676 4339 2682
rect 4345 2676 4348 2682
rect 4354 2676 4357 2682
rect 4363 2676 4373 2682
rect 4235 2675 4373 2676
rect 4235 2670 4243 2675
rect 4235 2664 4236 2670
rect 4242 2664 4243 2670
rect 4235 2661 4243 2664
rect 4235 2655 4236 2661
rect 4242 2655 4243 2661
rect 4235 2652 4243 2655
rect 4235 2646 4236 2652
rect 4242 2646 4243 2652
rect 4235 2636 4243 2646
rect 4679 2735 4687 2738
rect 4679 2729 4680 2735
rect 4686 2729 4687 2735
rect 4679 2726 4687 2729
rect 4679 2720 4680 2726
rect 4686 2720 4687 2726
rect 4679 2717 4687 2720
rect 4679 2711 4680 2717
rect 4686 2711 4687 2717
rect 4679 2708 4687 2711
rect 4679 2702 4680 2708
rect 4686 2702 4687 2708
rect 4679 2699 4687 2702
rect 4679 2693 4680 2699
rect 4686 2693 4687 2699
rect 4679 2690 4687 2693
rect 4679 2684 4680 2690
rect 4686 2684 4687 2690
rect 4679 2681 4687 2684
rect 4679 2675 4680 2681
rect 4686 2675 4687 2681
rect 4679 2672 4687 2675
rect 4679 2666 4680 2672
rect 4686 2666 4687 2672
rect 4679 2663 4687 2666
rect 4679 2657 4680 2663
rect 4686 2657 4687 2663
rect 4679 2654 4687 2657
rect 4679 2648 4680 2654
rect 4686 2648 4687 2654
rect 4679 2639 4687 2648
rect 6424 2792 6746 2793
rect 6424 2786 6434 2792
rect 6440 2786 6443 2792
rect 6449 2786 6452 2792
rect 6458 2786 6461 2792
rect 6467 2786 6472 2792
rect 6478 2786 6481 2792
rect 6487 2786 6490 2792
rect 6496 2786 6499 2792
rect 6505 2786 6508 2792
rect 6514 2786 6519 2792
rect 6525 2786 6528 2792
rect 6534 2786 6537 2792
rect 6543 2786 6546 2792
rect 6552 2786 6555 2792
rect 6561 2786 6564 2792
rect 6570 2786 6573 2792
rect 6579 2786 6582 2792
rect 6588 2786 6591 2792
rect 6597 2786 6602 2792
rect 6608 2786 6611 2792
rect 6617 2786 6620 2792
rect 6626 2786 6629 2792
rect 6635 2786 6638 2792
rect 6644 2786 6649 2792
rect 6655 2786 6658 2792
rect 6664 2786 6667 2792
rect 6673 2786 6676 2792
rect 6682 2786 6685 2792
rect 6691 2786 6694 2792
rect 6700 2786 6703 2792
rect 6709 2786 6712 2792
rect 6718 2786 6721 2792
rect 6727 2786 6730 2792
rect 6736 2786 6746 2792
rect 6424 2785 6746 2786
rect 6424 2783 6432 2785
rect 6424 2777 6425 2783
rect 6431 2777 6432 2783
rect 6424 2774 6432 2777
rect 6424 2768 6425 2774
rect 6431 2768 6432 2774
rect 6424 2765 6432 2768
rect 6424 2759 6425 2765
rect 6431 2759 6432 2765
rect 6738 2783 6746 2785
rect 6738 2777 6739 2783
rect 6745 2777 6746 2783
rect 6738 2774 6746 2777
rect 6738 2768 6739 2774
rect 6745 2768 6746 2774
rect 6738 2765 6746 2768
rect 6424 2756 6432 2759
rect 6738 2759 6739 2765
rect 6745 2759 6746 2765
rect 6424 2750 6425 2756
rect 6431 2750 6432 2756
rect 6424 2748 6432 2750
rect 6424 2742 6425 2748
rect 6431 2742 6432 2748
rect 6424 2739 6432 2742
rect 6424 2733 6425 2739
rect 6431 2733 6432 2739
rect 6424 2730 6432 2733
rect 6424 2724 6425 2730
rect 6431 2724 6432 2730
rect 6424 2721 6432 2724
rect 6424 2715 6425 2721
rect 6431 2715 6432 2721
rect 6424 2712 6432 2715
rect 6424 2706 6425 2712
rect 6431 2706 6432 2712
rect 6424 2704 6432 2706
rect 6294 2703 6432 2704
rect 6294 2697 6304 2703
rect 6310 2697 6313 2703
rect 6319 2697 6322 2703
rect 6328 2697 6331 2703
rect 6337 2697 6342 2703
rect 6348 2697 6351 2703
rect 6357 2697 6360 2703
rect 6366 2697 6369 2703
rect 6375 2697 6378 2703
rect 6384 2697 6389 2703
rect 6395 2697 6398 2703
rect 6404 2697 6407 2703
rect 6413 2697 6416 2703
rect 6422 2697 6432 2703
rect 6294 2696 6432 2697
rect 6294 2691 6302 2696
rect 6294 2685 6295 2691
rect 6301 2685 6302 2691
rect 6294 2682 6302 2685
rect 6294 2676 6295 2682
rect 6301 2676 6302 2682
rect 6294 2673 6302 2676
rect 6294 2667 6295 2673
rect 6301 2667 6302 2673
rect 6294 2657 6302 2667
rect 6738 2756 6746 2759
rect 6738 2750 6739 2756
rect 6745 2750 6746 2756
rect 6738 2747 6746 2750
rect 6738 2741 6739 2747
rect 6745 2741 6746 2747
rect 6738 2738 6746 2741
rect 6738 2732 6739 2738
rect 6745 2732 6746 2738
rect 6738 2729 6746 2732
rect 6738 2723 6739 2729
rect 6745 2723 6746 2729
rect 6738 2720 6746 2723
rect 6738 2714 6739 2720
rect 6745 2714 6746 2720
rect 6738 2711 6746 2714
rect 6738 2705 6739 2711
rect 6745 2705 6746 2711
rect 6738 2702 6746 2705
rect 6738 2696 6739 2702
rect 6745 2696 6746 2702
rect 6738 2693 6746 2696
rect 6738 2687 6739 2693
rect 6745 2687 6746 2693
rect 6738 2684 6746 2687
rect 6738 2678 6739 2684
rect 6745 2678 6746 2684
rect 6738 2675 6746 2678
rect 6738 2669 6739 2675
rect 6745 2669 6746 2675
rect 6738 2660 6746 2669
rect 8353 2774 8372 2797
rect 8353 2484 8372 2509
rect 3069 1910 3088 1935
rect 3069 1622 3088 1645
rect 8353 1928 8372 1951
rect 8353 1638 8372 1663
rect 3069 970 3088 995
rect 3069 682 3088 705
rect 4493 1022 4501 1031
rect 4493 1016 4494 1022
rect 4500 1016 4501 1022
rect 4493 1013 4501 1016
rect 4493 1007 4494 1013
rect 4500 1007 4501 1013
rect 4493 1004 4501 1007
rect 4493 998 4494 1004
rect 4500 998 4501 1004
rect 4493 995 4501 998
rect 4493 989 4494 995
rect 4500 989 4501 995
rect 4493 986 4501 989
rect 4493 980 4494 986
rect 4500 980 4501 986
rect 4493 977 4501 980
rect 4493 971 4494 977
rect 4500 971 4501 977
rect 4493 968 4501 971
rect 4493 962 4494 968
rect 4500 962 4501 968
rect 4493 959 4501 962
rect 4493 953 4494 959
rect 4500 953 4501 959
rect 4493 950 4501 953
rect 4493 944 4494 950
rect 4500 944 4501 950
rect 4493 941 4501 944
rect 4493 935 4494 941
rect 4500 935 4501 941
rect 4493 932 4501 935
rect 4937 1024 4945 1034
rect 4937 1018 4938 1024
rect 4944 1018 4945 1024
rect 4937 1015 4945 1018
rect 4937 1009 4938 1015
rect 4944 1009 4945 1015
rect 4937 1006 4945 1009
rect 4937 1000 4938 1006
rect 4944 1000 4945 1006
rect 4937 995 4945 1000
rect 4807 994 4945 995
rect 4807 988 4817 994
rect 4823 988 4826 994
rect 4832 988 4835 994
rect 4841 988 4844 994
rect 4850 988 4855 994
rect 4861 988 4864 994
rect 4870 988 4873 994
rect 4879 988 4882 994
rect 4888 988 4891 994
rect 4897 988 4902 994
rect 4908 988 4911 994
rect 4917 988 4920 994
rect 4926 988 4929 994
rect 4935 988 4945 994
rect 4807 987 4945 988
rect 4807 985 4815 987
rect 4807 979 4808 985
rect 4814 979 4815 985
rect 4807 976 4815 979
rect 4807 970 4808 976
rect 4814 970 4815 976
rect 4807 967 4815 970
rect 4807 961 4808 967
rect 4814 961 4815 967
rect 4807 958 4815 961
rect 4807 952 4808 958
rect 4814 952 4815 958
rect 4807 949 4815 952
rect 4807 943 4808 949
rect 4814 943 4815 949
rect 4807 941 4815 943
rect 4807 935 4808 941
rect 4814 935 4815 941
rect 4493 926 4494 932
rect 4500 926 4501 932
rect 4807 932 4815 935
rect 4493 923 4501 926
rect 4493 917 4494 923
rect 4500 917 4501 923
rect 4493 914 4501 917
rect 4493 908 4494 914
rect 4500 908 4501 914
rect 4493 906 4501 908
rect 4807 926 4808 932
rect 4814 926 4815 932
rect 4807 923 4815 926
rect 4807 917 4808 923
rect 4814 917 4815 923
rect 4807 914 4815 917
rect 4807 908 4808 914
rect 4814 908 4815 914
rect 4807 906 4815 908
rect 4493 905 4815 906
rect 4493 899 4503 905
rect 4509 899 4512 905
rect 4518 899 4521 905
rect 4527 899 4530 905
rect 4536 899 4539 905
rect 4545 899 4548 905
rect 4554 899 4557 905
rect 4563 899 4566 905
rect 4572 899 4575 905
rect 4581 899 4584 905
rect 4590 899 4595 905
rect 4601 899 4604 905
rect 4610 899 4613 905
rect 4619 899 4622 905
rect 4628 899 4631 905
rect 4637 899 4642 905
rect 4648 899 4651 905
rect 4657 899 4660 905
rect 4666 899 4669 905
rect 4675 899 4678 905
rect 4684 899 4687 905
rect 4693 899 4696 905
rect 4702 899 4705 905
rect 4711 899 4714 905
rect 4720 899 4725 905
rect 4731 899 4734 905
rect 4740 899 4743 905
rect 4749 899 4752 905
rect 4758 899 4761 905
rect 4767 899 4772 905
rect 4778 899 4781 905
rect 4787 899 4790 905
rect 4796 899 4799 905
rect 4805 899 4808 905
rect 4814 899 4815 905
rect 4493 898 4815 899
rect 6542 994 6550 1003
rect 6542 988 6543 994
rect 6549 988 6550 994
rect 6542 985 6550 988
rect 6542 979 6543 985
rect 6549 979 6550 985
rect 6542 976 6550 979
rect 6542 970 6543 976
rect 6549 970 6550 976
rect 6542 967 6550 970
rect 6542 961 6543 967
rect 6549 961 6550 967
rect 6542 958 6550 961
rect 6542 952 6543 958
rect 6549 952 6550 958
rect 6542 949 6550 952
rect 6542 943 6543 949
rect 6549 943 6550 949
rect 6542 940 6550 943
rect 6542 934 6543 940
rect 6549 934 6550 940
rect 6542 931 6550 934
rect 6542 925 6543 931
rect 6549 925 6550 931
rect 6542 922 6550 925
rect 6542 916 6543 922
rect 6549 916 6550 922
rect 6542 913 6550 916
rect 6542 907 6543 913
rect 6549 907 6550 913
rect 6542 904 6550 907
rect 6986 996 6994 1006
rect 6986 990 6987 996
rect 6993 990 6994 996
rect 6986 987 6994 990
rect 6986 981 6987 987
rect 6993 981 6994 987
rect 6986 978 6994 981
rect 6986 972 6987 978
rect 6993 972 6994 978
rect 6986 967 6994 972
rect 6856 966 6994 967
rect 6856 960 6866 966
rect 6872 960 6875 966
rect 6881 960 6884 966
rect 6890 960 6893 966
rect 6899 960 6904 966
rect 6910 960 6913 966
rect 6919 960 6922 966
rect 6928 960 6931 966
rect 6937 960 6940 966
rect 6946 960 6951 966
rect 6957 960 6960 966
rect 6966 960 6969 966
rect 6975 960 6978 966
rect 6984 960 6994 966
rect 6856 959 6994 960
rect 6856 957 6864 959
rect 6856 951 6857 957
rect 6863 951 6864 957
rect 6856 948 6864 951
rect 6856 942 6857 948
rect 6863 942 6864 948
rect 6856 939 6864 942
rect 6856 933 6857 939
rect 6863 933 6864 939
rect 6856 930 6864 933
rect 6856 924 6857 930
rect 6863 924 6864 930
rect 6856 921 6864 924
rect 6856 915 6857 921
rect 6863 915 6864 921
rect 6856 913 6864 915
rect 6856 907 6857 913
rect 6863 907 6864 913
rect 6542 898 6543 904
rect 6549 898 6550 904
rect 6856 904 6864 907
rect 6542 895 6550 898
rect 6542 889 6543 895
rect 6549 889 6550 895
rect 6542 886 6550 889
rect 6542 880 6543 886
rect 6549 880 6550 886
rect 6542 878 6550 880
rect 6856 898 6857 904
rect 6863 898 6864 904
rect 6856 895 6864 898
rect 6856 889 6857 895
rect 6863 889 6864 895
rect 6856 886 6864 889
rect 6856 880 6857 886
rect 6863 880 6864 886
rect 6856 878 6864 880
rect 6542 877 6864 878
rect 6542 871 6552 877
rect 6558 871 6561 877
rect 6567 871 6570 877
rect 6576 871 6579 877
rect 6585 871 6588 877
rect 6594 871 6597 877
rect 6603 871 6606 877
rect 6612 871 6615 877
rect 6621 871 6624 877
rect 6630 871 6633 877
rect 6639 871 6644 877
rect 6650 871 6653 877
rect 6659 871 6662 877
rect 6668 871 6671 877
rect 6677 871 6680 877
rect 6686 871 6691 877
rect 6697 871 6700 877
rect 6706 871 6709 877
rect 6715 871 6718 877
rect 6724 871 6727 877
rect 6733 871 6736 877
rect 6742 871 6745 877
rect 6751 871 6754 877
rect 6760 871 6763 877
rect 6769 871 6774 877
rect 6780 871 6783 877
rect 6789 871 6792 877
rect 6798 871 6801 877
rect 6807 871 6810 877
rect 6816 871 6821 877
rect 6827 871 6830 877
rect 6836 871 6839 877
rect 6845 871 6848 877
rect 6854 871 6864 877
rect 6542 870 6864 871
rect 8352 924 8371 947
rect 8352 634 8371 659
rect 3917 -391 3942 -372
rect 4207 -391 4230 -372
rect 5071 -390 5096 -371
rect 5361 -390 5384 -371
rect 6222 -390 6247 -371
rect 6512 -390 6535 -371
rect 7313 -390 7338 -371
rect 7603 -390 7626 -371
<< psubstratepcontact >>
rect 3887 3436 3909 3585
rect 3928 3436 4203 3457
rect 4222 3436 4244 3585
rect 5052 3436 5074 3585
rect 5093 3436 5368 3457
rect 5387 3436 5409 3585
rect 6207 3436 6229 3585
rect 6248 3436 6523 3457
rect 6542 3436 6564 3585
rect 7400 3436 7422 3585
rect 7441 3436 7716 3457
rect 7735 3436 7757 3585
rect 3335 2847 3484 2869
rect 3463 2553 3484 2828
rect 6415 2800 6421 2806
rect 6424 2800 6430 2806
rect 4356 2779 4362 2785
rect 4365 2779 4371 2785
rect 4446 2779 4452 2785
rect 4455 2779 4461 2785
rect 4464 2779 4470 2785
rect 4473 2779 4479 2785
rect 4482 2779 4488 2785
rect 4491 2779 4497 2785
rect 4500 2779 4506 2785
rect 4509 2779 4515 2785
rect 4518 2779 4524 2785
rect 4527 2779 4533 2785
rect 4536 2779 4542 2785
rect 4545 2779 4551 2785
rect 4554 2779 4560 2785
rect 4563 2779 4569 2785
rect 4572 2779 4578 2785
rect 4581 2779 4587 2785
rect 4590 2779 4596 2785
rect 4599 2779 4605 2785
rect 4608 2779 4614 2785
rect 4617 2779 4623 2785
rect 4626 2779 4632 2785
rect 4635 2779 4641 2785
rect 4644 2779 4650 2785
rect 4653 2779 4659 2785
rect 4662 2779 4668 2785
rect 4671 2779 4677 2785
rect 4680 2779 4686 2785
rect 4689 2779 4695 2785
rect 4347 2770 4353 2776
rect 4347 2761 4353 2767
rect 4347 2752 4353 2758
rect 4347 2743 4353 2749
rect 4347 2735 4353 2741
rect 4347 2726 4353 2732
rect 4347 2717 4353 2723
rect 4347 2708 4353 2714
rect 4347 2699 4353 2705
rect 4231 2690 4237 2696
rect 4240 2690 4246 2696
rect 4249 2690 4255 2696
rect 4258 2690 4264 2696
rect 4267 2690 4273 2696
rect 4276 2690 4282 2696
rect 4285 2690 4291 2696
rect 4294 2690 4300 2696
rect 4303 2690 4309 2696
rect 4312 2690 4318 2696
rect 4321 2690 4327 2696
rect 4330 2690 4336 2696
rect 4339 2690 4345 2696
rect 4222 2682 4228 2688
rect 4222 2673 4228 2679
rect 4222 2664 4228 2670
rect 4222 2655 4228 2661
rect 4222 2646 4228 2652
rect 4698 2770 4704 2776
rect 4698 2761 4704 2767
rect 4698 2752 4704 2758
rect 4698 2743 4704 2749
rect 4698 2731 4704 2737
rect 4698 2722 4704 2728
rect 4698 2713 4704 2719
rect 4698 2704 4704 2710
rect 4698 2697 4704 2703
rect 4698 2688 4704 2694
rect 4698 2679 4704 2685
rect 4698 2670 4704 2676
rect 4698 2661 4704 2667
rect 4698 2652 4704 2658
rect 6505 2800 6511 2806
rect 6514 2800 6520 2806
rect 6523 2800 6529 2806
rect 6532 2800 6538 2806
rect 6541 2800 6547 2806
rect 6550 2800 6556 2806
rect 6559 2800 6565 2806
rect 6568 2800 6574 2806
rect 6577 2800 6583 2806
rect 6586 2800 6592 2806
rect 6595 2800 6601 2806
rect 6604 2800 6610 2806
rect 6613 2800 6619 2806
rect 6622 2800 6628 2806
rect 6631 2800 6637 2806
rect 6640 2800 6646 2806
rect 6649 2800 6655 2806
rect 6658 2800 6664 2806
rect 6667 2800 6673 2806
rect 6676 2800 6682 2806
rect 6685 2800 6691 2806
rect 6694 2800 6700 2806
rect 6703 2800 6709 2806
rect 6712 2800 6718 2806
rect 6721 2800 6727 2806
rect 6730 2800 6736 2806
rect 6739 2800 6745 2806
rect 6748 2800 6754 2806
rect 6406 2791 6412 2797
rect 6406 2782 6412 2788
rect 6406 2773 6412 2779
rect 6406 2764 6412 2770
rect 6406 2756 6412 2762
rect 6406 2747 6412 2753
rect 6406 2738 6412 2744
rect 6406 2729 6412 2735
rect 6406 2720 6412 2726
rect 6290 2711 6296 2717
rect 6299 2711 6305 2717
rect 6308 2711 6314 2717
rect 6317 2711 6323 2717
rect 6326 2711 6332 2717
rect 6335 2711 6341 2717
rect 6344 2711 6350 2717
rect 6353 2711 6359 2717
rect 6362 2711 6368 2717
rect 6371 2711 6377 2717
rect 6380 2711 6386 2717
rect 6389 2711 6395 2717
rect 6398 2711 6404 2717
rect 6281 2703 6287 2709
rect 6281 2694 6287 2700
rect 6281 2685 6287 2691
rect 6281 2676 6287 2682
rect 6281 2667 6287 2673
rect 4222 2583 4228 2589
rect 4231 2575 4237 2581
rect 4240 2575 4246 2581
rect 4249 2575 4255 2581
rect 4258 2575 4264 2581
rect 4267 2575 4273 2581
rect 4276 2575 4282 2581
rect 4285 2575 4291 2581
rect 4294 2575 4300 2581
rect 4303 2575 4309 2581
rect 4312 2575 4318 2581
rect 4321 2575 4327 2581
rect 4330 2575 4336 2581
rect 4339 2575 4345 2581
rect 4348 2575 4354 2581
rect 4355 2575 4361 2581
rect 4362 2566 4368 2572
rect 4362 2557 4368 2563
rect 4371 2550 4377 2556
rect 4380 2550 4386 2556
rect 4389 2550 4395 2556
rect 4398 2550 4404 2556
rect 4407 2550 4413 2556
rect 4416 2550 4422 2556
rect 4425 2550 4431 2556
rect 4434 2550 4440 2556
rect 4443 2550 4449 2556
rect 4452 2550 4458 2556
rect 4461 2550 4467 2556
rect 3335 2512 3484 2534
rect 4468 2541 4474 2547
rect 4468 2532 4474 2538
rect 4468 2523 4474 2529
rect 4468 2514 4474 2520
rect 4609 2608 4615 2614
rect 4618 2608 4624 2614
rect 4627 2608 4633 2614
rect 4636 2608 4642 2614
rect 4645 2608 4651 2614
rect 4654 2608 4660 2614
rect 4663 2608 4669 2614
rect 4672 2608 4678 2614
rect 4681 2608 4687 2614
rect 4690 2608 4696 2614
rect 6757 2791 6763 2797
rect 6757 2782 6763 2788
rect 6757 2773 6763 2779
rect 6757 2764 6763 2770
rect 6757 2752 6763 2758
rect 6757 2743 6763 2749
rect 6757 2734 6763 2740
rect 6757 2725 6763 2731
rect 6757 2718 6763 2724
rect 6757 2709 6763 2715
rect 6757 2700 6763 2706
rect 6757 2691 6763 2697
rect 6757 2682 6763 2688
rect 6757 2673 6763 2679
rect 4600 2599 4606 2605
rect 4600 2590 4606 2596
rect 6281 2604 6287 2610
rect 6290 2596 6296 2602
rect 6299 2596 6305 2602
rect 6308 2596 6314 2602
rect 6317 2596 6323 2602
rect 6326 2596 6332 2602
rect 6335 2596 6341 2602
rect 6344 2596 6350 2602
rect 6353 2596 6359 2602
rect 6362 2596 6368 2602
rect 6371 2596 6377 2602
rect 6380 2596 6386 2602
rect 6389 2596 6395 2602
rect 6398 2596 6404 2602
rect 6407 2596 6413 2602
rect 6414 2596 6420 2602
rect 4600 2581 4606 2587
rect 4600 2572 4606 2578
rect 6421 2587 6427 2593
rect 6421 2578 6427 2584
rect 6430 2571 6436 2577
rect 6439 2571 6445 2577
rect 6448 2571 6454 2577
rect 6457 2571 6463 2577
rect 6466 2571 6472 2577
rect 6475 2571 6481 2577
rect 6484 2571 6490 2577
rect 6493 2571 6499 2577
rect 6502 2571 6508 2577
rect 6511 2571 6517 2577
rect 6520 2571 6526 2577
rect 4600 2563 4606 2569
rect 4600 2554 4606 2560
rect 4600 2545 4606 2551
rect 4600 2536 4606 2542
rect 4600 2527 4606 2533
rect 4600 2518 4606 2524
rect 4468 2505 4474 2511
rect 4468 2496 4474 2502
rect 4600 2509 4606 2515
rect 4600 2500 4606 2506
rect 6527 2562 6533 2568
rect 6527 2553 6533 2559
rect 6527 2544 6533 2550
rect 6527 2535 6533 2541
rect 6668 2629 6674 2635
rect 6677 2629 6683 2635
rect 6686 2629 6692 2635
rect 6695 2629 6701 2635
rect 6704 2629 6710 2635
rect 6713 2629 6719 2635
rect 6722 2629 6728 2635
rect 6731 2629 6737 2635
rect 6740 2629 6746 2635
rect 6749 2629 6755 2635
rect 7958 2795 8107 2817
rect 6659 2620 6665 2626
rect 6659 2611 6665 2617
rect 6659 2602 6665 2608
rect 6659 2593 6665 2599
rect 6659 2584 6665 2590
rect 6659 2575 6665 2581
rect 6659 2566 6665 2572
rect 6659 2557 6665 2563
rect 6659 2548 6665 2554
rect 6659 2539 6665 2545
rect 6527 2526 6533 2532
rect 6527 2517 6533 2523
rect 6659 2530 6665 2536
rect 6659 2521 6665 2527
rect 6659 2512 6665 2518
rect 6536 2505 6542 2511
rect 6545 2505 6551 2511
rect 6554 2505 6560 2511
rect 6563 2505 6569 2511
rect 6572 2505 6578 2511
rect 6581 2505 6587 2511
rect 6590 2505 6596 2511
rect 6599 2505 6605 2511
rect 6608 2505 6614 2511
rect 6617 2505 6623 2511
rect 6626 2505 6632 2511
rect 6635 2505 6641 2511
rect 6644 2505 6650 2511
rect 6653 2505 6659 2511
rect 4600 2491 4606 2497
rect 7958 2501 7979 2776
rect 4477 2484 4483 2490
rect 4486 2484 4492 2490
rect 4495 2484 4501 2490
rect 4504 2484 4510 2490
rect 4513 2484 4519 2490
rect 4522 2484 4528 2490
rect 4531 2484 4537 2490
rect 4540 2484 4546 2490
rect 4549 2484 4555 2490
rect 4558 2484 4564 2490
rect 4567 2484 4573 2490
rect 4576 2484 4582 2490
rect 4585 2484 4591 2490
rect 4594 2484 4600 2490
rect 7958 2460 8107 2482
rect 3334 1937 3483 1959
rect 3462 1643 3483 1918
rect 3334 1602 3483 1624
rect 7958 1949 8107 1971
rect 7958 1655 7979 1930
rect 7958 1614 8107 1636
rect 4580 1180 4586 1186
rect 4589 1180 4595 1186
rect 4598 1180 4604 1186
rect 4607 1180 4613 1186
rect 4616 1180 4622 1186
rect 4625 1180 4631 1186
rect 4634 1180 4640 1186
rect 4643 1180 4649 1186
rect 4652 1180 4658 1186
rect 4661 1180 4667 1186
rect 4670 1180 4676 1186
rect 4679 1180 4685 1186
rect 4688 1180 4694 1186
rect 4697 1180 4703 1186
rect 4574 1173 4580 1179
rect 4574 1164 4580 1170
rect 4574 1155 4580 1161
rect 4706 1168 4712 1174
rect 4706 1159 4712 1165
rect 4574 1146 4580 1152
rect 4574 1137 4580 1143
rect 4574 1128 4580 1134
rect 4574 1119 4580 1125
rect 4574 1110 4580 1116
rect 4574 1101 4580 1107
rect 4574 1092 4580 1098
rect 4574 1083 4580 1089
rect 4574 1074 4580 1080
rect 4574 1065 4580 1071
rect 4484 1056 4490 1062
rect 4493 1056 4499 1062
rect 4502 1056 4508 1062
rect 4511 1056 4517 1062
rect 4520 1056 4526 1062
rect 4529 1056 4535 1062
rect 4538 1056 4544 1062
rect 4547 1056 4553 1062
rect 4556 1056 4562 1062
rect 4565 1056 4571 1062
rect 4706 1150 4712 1156
rect 4706 1141 4712 1147
rect 4706 1132 4712 1138
rect 4706 1123 4712 1129
rect 6629 1152 6635 1158
rect 6638 1152 6644 1158
rect 6647 1152 6653 1158
rect 6656 1152 6662 1158
rect 6665 1152 6671 1158
rect 6674 1152 6680 1158
rect 6683 1152 6689 1158
rect 6692 1152 6698 1158
rect 6701 1152 6707 1158
rect 6710 1152 6716 1158
rect 6719 1152 6725 1158
rect 6728 1152 6734 1158
rect 6737 1152 6743 1158
rect 6746 1152 6752 1158
rect 6623 1145 6629 1151
rect 6623 1136 6629 1142
rect 6623 1127 6629 1133
rect 6755 1140 6761 1146
rect 6755 1131 6761 1137
rect 4713 1114 4719 1120
rect 4722 1114 4728 1120
rect 4731 1114 4737 1120
rect 4740 1114 4746 1120
rect 4749 1114 4755 1120
rect 4758 1114 4764 1120
rect 4767 1114 4773 1120
rect 4776 1114 4782 1120
rect 4785 1114 4791 1120
rect 4794 1114 4800 1120
rect 4803 1114 4809 1120
rect 4812 1107 4818 1113
rect 4812 1098 4818 1104
rect 6623 1118 6629 1124
rect 6623 1109 6629 1115
rect 6623 1100 6629 1106
rect 4819 1089 4825 1095
rect 4826 1089 4832 1095
rect 4835 1089 4841 1095
rect 4844 1089 4850 1095
rect 4853 1089 4859 1095
rect 4862 1089 4868 1095
rect 4871 1089 4877 1095
rect 4880 1089 4886 1095
rect 4889 1089 4895 1095
rect 4898 1089 4904 1095
rect 4907 1089 4913 1095
rect 4916 1089 4922 1095
rect 4925 1089 4931 1095
rect 4934 1089 4940 1095
rect 4943 1089 4949 1095
rect 4952 1081 4958 1087
rect 3334 997 3483 1019
rect 3462 703 3483 978
rect 4476 1012 4482 1018
rect 4476 1003 4482 1009
rect 4476 994 4482 1000
rect 4476 985 4482 991
rect 4476 976 4482 982
rect 4476 967 4482 973
rect 4476 960 4482 966
rect 4476 951 4482 957
rect 4476 942 4482 948
rect 4476 933 4482 939
rect 4476 921 4482 927
rect 4476 912 4482 918
rect 4476 903 4482 909
rect 4476 894 4482 900
rect 6623 1091 6629 1097
rect 6623 1082 6629 1088
rect 6623 1073 6629 1079
rect 6623 1064 6629 1070
rect 6623 1055 6629 1061
rect 6623 1046 6629 1052
rect 6623 1037 6629 1043
rect 4952 1018 4958 1024
rect 4952 1009 4958 1015
rect 4952 1000 4958 1006
rect 4952 991 4958 997
rect 4952 982 4958 988
rect 4835 974 4841 980
rect 4844 974 4850 980
rect 4853 974 4859 980
rect 4862 974 4868 980
rect 4871 974 4877 980
rect 4880 974 4886 980
rect 4889 974 4895 980
rect 4898 974 4904 980
rect 4907 974 4913 980
rect 4916 974 4922 980
rect 4925 974 4931 980
rect 4934 974 4940 980
rect 4943 974 4949 980
rect 6533 1028 6539 1034
rect 6542 1028 6548 1034
rect 6551 1028 6557 1034
rect 6560 1028 6566 1034
rect 6569 1028 6575 1034
rect 6578 1028 6584 1034
rect 6587 1028 6593 1034
rect 6596 1028 6602 1034
rect 6605 1028 6611 1034
rect 6614 1028 6620 1034
rect 6755 1122 6761 1128
rect 6755 1113 6761 1119
rect 6755 1104 6761 1110
rect 6755 1095 6761 1101
rect 6762 1086 6768 1092
rect 6771 1086 6777 1092
rect 6780 1086 6786 1092
rect 6789 1086 6795 1092
rect 6798 1086 6804 1092
rect 6807 1086 6813 1092
rect 6816 1086 6822 1092
rect 6825 1086 6831 1092
rect 6834 1086 6840 1092
rect 6843 1086 6849 1092
rect 6852 1086 6858 1092
rect 6861 1079 6867 1085
rect 6861 1070 6867 1076
rect 6868 1061 6874 1067
rect 6875 1061 6881 1067
rect 6884 1061 6890 1067
rect 6893 1061 6899 1067
rect 6902 1061 6908 1067
rect 6911 1061 6917 1067
rect 6920 1061 6926 1067
rect 6929 1061 6935 1067
rect 6938 1061 6944 1067
rect 6947 1061 6953 1067
rect 6956 1061 6962 1067
rect 6965 1061 6971 1067
rect 6974 1061 6980 1067
rect 6983 1061 6989 1067
rect 6992 1061 6998 1067
rect 7001 1053 7007 1059
rect 6525 984 6531 990
rect 6525 975 6531 981
rect 4827 965 4833 971
rect 4827 956 4833 962
rect 4827 947 4833 953
rect 4827 938 4833 944
rect 4827 929 4833 935
rect 4827 921 4833 927
rect 4827 912 4833 918
rect 4827 903 4833 909
rect 4827 894 4833 900
rect 4485 885 4491 891
rect 4494 885 4500 891
rect 4503 885 4509 891
rect 4512 885 4518 891
rect 4521 885 4527 891
rect 4530 885 4536 891
rect 4539 885 4545 891
rect 4548 885 4554 891
rect 4557 885 4563 891
rect 4566 885 4572 891
rect 4575 885 4581 891
rect 4584 885 4590 891
rect 4593 885 4599 891
rect 4602 885 4608 891
rect 4611 885 4617 891
rect 4620 885 4626 891
rect 4629 885 4635 891
rect 4638 885 4644 891
rect 4647 885 4653 891
rect 4656 885 4662 891
rect 4665 885 4671 891
rect 4674 885 4680 891
rect 4683 885 4689 891
rect 4692 885 4698 891
rect 4701 885 4707 891
rect 4710 885 4716 891
rect 4719 885 4725 891
rect 4728 885 4734 891
rect 4809 885 4815 891
rect 4818 885 4824 891
rect 6525 966 6531 972
rect 6525 957 6531 963
rect 6525 948 6531 954
rect 6525 939 6531 945
rect 6525 932 6531 938
rect 6525 923 6531 929
rect 6525 914 6531 920
rect 6525 905 6531 911
rect 6525 893 6531 899
rect 6525 884 6531 890
rect 6525 875 6531 881
rect 6525 866 6531 872
rect 7001 990 7007 996
rect 7001 981 7007 987
rect 7001 972 7007 978
rect 7001 963 7007 969
rect 7001 954 7007 960
rect 6884 946 6890 952
rect 6893 946 6899 952
rect 6902 946 6908 952
rect 6911 946 6917 952
rect 6920 946 6926 952
rect 6929 946 6935 952
rect 6938 946 6944 952
rect 6947 946 6953 952
rect 6956 946 6962 952
rect 6965 946 6971 952
rect 6974 946 6980 952
rect 6983 946 6989 952
rect 6992 946 6998 952
rect 7957 945 8106 967
rect 6876 937 6882 943
rect 6876 928 6882 934
rect 6876 919 6882 925
rect 6876 910 6882 916
rect 6876 901 6882 907
rect 6876 893 6882 899
rect 6876 884 6882 890
rect 6876 875 6882 881
rect 6876 866 6882 872
rect 6534 857 6540 863
rect 6543 857 6549 863
rect 6552 857 6558 863
rect 6561 857 6567 863
rect 6570 857 6576 863
rect 6579 857 6585 863
rect 6588 857 6594 863
rect 6597 857 6603 863
rect 6606 857 6612 863
rect 6615 857 6621 863
rect 6624 857 6630 863
rect 6633 857 6639 863
rect 6642 857 6648 863
rect 6651 857 6657 863
rect 6660 857 6666 863
rect 6669 857 6675 863
rect 6678 857 6684 863
rect 6687 857 6693 863
rect 6696 857 6702 863
rect 6705 857 6711 863
rect 6714 857 6720 863
rect 6723 857 6729 863
rect 6732 857 6738 863
rect 6741 857 6747 863
rect 6750 857 6756 863
rect 6759 857 6765 863
rect 6768 857 6774 863
rect 6777 857 6783 863
rect 6849 857 6855 863
rect 6858 857 6864 863
rect 6867 857 6873 863
rect 3334 662 3483 684
rect 7957 651 7978 926
rect 7957 610 8106 632
rect 3893 -126 3915 23
rect 3934 2 4209 23
rect 4228 -126 4250 23
rect 5047 -125 5069 24
rect 5088 3 5363 24
rect 5382 -125 5404 24
rect 6198 -125 6220 24
rect 6239 3 6514 24
rect 6533 -125 6555 24
rect 7289 -125 7311 24
rect 7330 3 7605 24
rect 7624 -125 7646 24
<< nsubstratencontact >>
rect 3886 3701 3907 3850
rect 3930 3831 4195 3850
rect 4220 3701 4241 3850
rect 5051 3701 5072 3850
rect 5095 3831 5360 3850
rect 5385 3701 5406 3850
rect 6206 3701 6227 3850
rect 6250 3831 6515 3850
rect 6540 3701 6561 3850
rect 7399 3701 7420 3850
rect 7443 3831 7708 3850
rect 7733 3701 7754 3850
rect 3070 2845 3219 2866
rect 3070 2555 3089 2820
rect 4375 2765 4381 2771
rect 4384 2765 4390 2771
rect 4393 2765 4399 2771
rect 4402 2765 4408 2771
rect 4413 2765 4419 2771
rect 4422 2765 4428 2771
rect 4431 2765 4437 2771
rect 4440 2765 4446 2771
rect 4449 2765 4455 2771
rect 4460 2765 4466 2771
rect 4469 2765 4475 2771
rect 4478 2765 4484 2771
rect 4487 2765 4493 2771
rect 4496 2765 4502 2771
rect 4505 2765 4511 2771
rect 4514 2765 4520 2771
rect 4523 2765 4529 2771
rect 4532 2765 4538 2771
rect 4543 2765 4549 2771
rect 4552 2765 4558 2771
rect 4561 2765 4567 2771
rect 4570 2765 4576 2771
rect 4579 2765 4585 2771
rect 4590 2765 4596 2771
rect 4599 2765 4605 2771
rect 4608 2765 4614 2771
rect 4617 2765 4623 2771
rect 4626 2765 4632 2771
rect 4635 2765 4641 2771
rect 4644 2765 4650 2771
rect 4653 2765 4659 2771
rect 4662 2765 4668 2771
rect 4671 2765 4677 2771
rect 4366 2756 4372 2762
rect 4366 2747 4372 2753
rect 4366 2738 4372 2744
rect 4680 2756 4686 2762
rect 4680 2747 4686 2753
rect 4680 2738 4686 2744
rect 4366 2729 4372 2735
rect 4366 2721 4372 2727
rect 4366 2712 4372 2718
rect 4366 2703 4372 2709
rect 4366 2694 4372 2700
rect 4366 2685 4372 2691
rect 4245 2676 4251 2682
rect 4254 2676 4260 2682
rect 4263 2676 4269 2682
rect 4272 2676 4278 2682
rect 4283 2676 4289 2682
rect 4292 2676 4298 2682
rect 4301 2676 4307 2682
rect 4310 2676 4316 2682
rect 4319 2676 4325 2682
rect 4330 2676 4336 2682
rect 4339 2676 4345 2682
rect 4348 2676 4354 2682
rect 4357 2676 4363 2682
rect 4236 2664 4242 2670
rect 4236 2655 4242 2661
rect 4236 2646 4242 2652
rect 4680 2729 4686 2735
rect 4680 2720 4686 2726
rect 4680 2711 4686 2717
rect 4680 2702 4686 2708
rect 4680 2693 4686 2699
rect 4680 2684 4686 2690
rect 4680 2675 4686 2681
rect 4680 2666 4686 2672
rect 4680 2657 4686 2663
rect 4680 2648 4686 2654
rect 6434 2786 6440 2792
rect 6443 2786 6449 2792
rect 6452 2786 6458 2792
rect 6461 2786 6467 2792
rect 6472 2786 6478 2792
rect 6481 2786 6487 2792
rect 6490 2786 6496 2792
rect 6499 2786 6505 2792
rect 6508 2786 6514 2792
rect 6519 2786 6525 2792
rect 6528 2786 6534 2792
rect 6537 2786 6543 2792
rect 6546 2786 6552 2792
rect 6555 2786 6561 2792
rect 6564 2786 6570 2792
rect 6573 2786 6579 2792
rect 6582 2786 6588 2792
rect 6591 2786 6597 2792
rect 6602 2786 6608 2792
rect 6611 2786 6617 2792
rect 6620 2786 6626 2792
rect 6629 2786 6635 2792
rect 6638 2786 6644 2792
rect 6649 2786 6655 2792
rect 6658 2786 6664 2792
rect 6667 2786 6673 2792
rect 6676 2786 6682 2792
rect 6685 2786 6691 2792
rect 6694 2786 6700 2792
rect 6703 2786 6709 2792
rect 6712 2786 6718 2792
rect 6721 2786 6727 2792
rect 6730 2786 6736 2792
rect 6425 2777 6431 2783
rect 6425 2768 6431 2774
rect 6425 2759 6431 2765
rect 6739 2777 6745 2783
rect 6739 2768 6745 2774
rect 6739 2759 6745 2765
rect 6425 2750 6431 2756
rect 6425 2742 6431 2748
rect 6425 2733 6431 2739
rect 6425 2724 6431 2730
rect 6425 2715 6431 2721
rect 6425 2706 6431 2712
rect 3070 2511 3219 2532
rect 6304 2697 6310 2703
rect 6313 2697 6319 2703
rect 6322 2697 6328 2703
rect 6331 2697 6337 2703
rect 6342 2697 6348 2703
rect 6351 2697 6357 2703
rect 6360 2697 6366 2703
rect 6369 2697 6375 2703
rect 6378 2697 6384 2703
rect 6389 2697 6395 2703
rect 6398 2697 6404 2703
rect 6407 2697 6413 2703
rect 6416 2697 6422 2703
rect 6295 2685 6301 2691
rect 6295 2676 6301 2682
rect 6295 2667 6301 2673
rect 6739 2750 6745 2756
rect 6739 2741 6745 2747
rect 6739 2732 6745 2738
rect 6739 2723 6745 2729
rect 6739 2714 6745 2720
rect 6739 2705 6745 2711
rect 6739 2696 6745 2702
rect 6739 2687 6745 2693
rect 6739 2678 6745 2684
rect 6739 2669 6745 2675
rect 8223 2797 8372 2818
rect 8353 2509 8372 2774
rect 8223 2463 8372 2484
rect 3069 1935 3218 1956
rect 3069 1645 3088 1910
rect 3069 1601 3218 1622
rect 8223 1951 8372 1972
rect 8353 1663 8372 1928
rect 8223 1617 8372 1638
rect 3069 995 3218 1016
rect 3069 705 3088 970
rect 4494 1016 4500 1022
rect 4494 1007 4500 1013
rect 4494 998 4500 1004
rect 4494 989 4500 995
rect 4494 980 4500 986
rect 4494 971 4500 977
rect 4494 962 4500 968
rect 4494 953 4500 959
rect 4494 944 4500 950
rect 4494 935 4500 941
rect 4938 1018 4944 1024
rect 4938 1009 4944 1015
rect 4938 1000 4944 1006
rect 4817 988 4823 994
rect 4826 988 4832 994
rect 4835 988 4841 994
rect 4844 988 4850 994
rect 4855 988 4861 994
rect 4864 988 4870 994
rect 4873 988 4879 994
rect 4882 988 4888 994
rect 4891 988 4897 994
rect 4902 988 4908 994
rect 4911 988 4917 994
rect 4920 988 4926 994
rect 4929 988 4935 994
rect 4808 979 4814 985
rect 4808 970 4814 976
rect 4808 961 4814 967
rect 4808 952 4814 958
rect 4808 943 4814 949
rect 4808 935 4814 941
rect 4494 926 4500 932
rect 4494 917 4500 923
rect 4494 908 4500 914
rect 4808 926 4814 932
rect 4808 917 4814 923
rect 4808 908 4814 914
rect 4503 899 4509 905
rect 4512 899 4518 905
rect 4521 899 4527 905
rect 4530 899 4536 905
rect 4539 899 4545 905
rect 4548 899 4554 905
rect 4557 899 4563 905
rect 4566 899 4572 905
rect 4575 899 4581 905
rect 4584 899 4590 905
rect 4595 899 4601 905
rect 4604 899 4610 905
rect 4613 899 4619 905
rect 4622 899 4628 905
rect 4631 899 4637 905
rect 4642 899 4648 905
rect 4651 899 4657 905
rect 4660 899 4666 905
rect 4669 899 4675 905
rect 4678 899 4684 905
rect 4687 899 4693 905
rect 4696 899 4702 905
rect 4705 899 4711 905
rect 4714 899 4720 905
rect 4725 899 4731 905
rect 4734 899 4740 905
rect 4743 899 4749 905
rect 4752 899 4758 905
rect 4761 899 4767 905
rect 4772 899 4778 905
rect 4781 899 4787 905
rect 4790 899 4796 905
rect 4799 899 4805 905
rect 4808 899 4814 905
rect 6543 988 6549 994
rect 6543 979 6549 985
rect 6543 970 6549 976
rect 6543 961 6549 967
rect 6543 952 6549 958
rect 6543 943 6549 949
rect 6543 934 6549 940
rect 6543 925 6549 931
rect 6543 916 6549 922
rect 6543 907 6549 913
rect 6987 990 6993 996
rect 6987 981 6993 987
rect 6987 972 6993 978
rect 6866 960 6872 966
rect 6875 960 6881 966
rect 6884 960 6890 966
rect 6893 960 6899 966
rect 6904 960 6910 966
rect 6913 960 6919 966
rect 6922 960 6928 966
rect 6931 960 6937 966
rect 6940 960 6946 966
rect 6951 960 6957 966
rect 6960 960 6966 966
rect 6969 960 6975 966
rect 6978 960 6984 966
rect 6857 951 6863 957
rect 6857 942 6863 948
rect 6857 933 6863 939
rect 6857 924 6863 930
rect 6857 915 6863 921
rect 6857 907 6863 913
rect 6543 898 6549 904
rect 6543 889 6549 895
rect 6543 880 6549 886
rect 6857 898 6863 904
rect 6857 889 6863 895
rect 6857 880 6863 886
rect 6552 871 6558 877
rect 6561 871 6567 877
rect 6570 871 6576 877
rect 6579 871 6585 877
rect 6588 871 6594 877
rect 6597 871 6603 877
rect 6606 871 6612 877
rect 6615 871 6621 877
rect 6624 871 6630 877
rect 6633 871 6639 877
rect 6644 871 6650 877
rect 6653 871 6659 877
rect 6662 871 6668 877
rect 6671 871 6677 877
rect 6680 871 6686 877
rect 6691 871 6697 877
rect 6700 871 6706 877
rect 6709 871 6715 877
rect 6718 871 6724 877
rect 6727 871 6733 877
rect 6736 871 6742 877
rect 6745 871 6751 877
rect 6754 871 6760 877
rect 6763 871 6769 877
rect 6774 871 6780 877
rect 6783 871 6789 877
rect 6792 871 6798 877
rect 6801 871 6807 877
rect 6810 871 6816 877
rect 6821 871 6827 877
rect 6830 871 6836 877
rect 6839 871 6845 877
rect 6848 871 6854 877
rect 8222 947 8371 968
rect 3069 661 3218 682
rect 8352 659 8371 924
rect 8222 613 8371 634
rect 3896 -391 3917 -242
rect 3942 -391 4207 -372
rect 4230 -391 4251 -242
rect 5050 -390 5071 -241
rect 5096 -390 5361 -371
rect 5384 -390 5405 -241
rect 6201 -390 6222 -241
rect 6247 -390 6512 -371
rect 6535 -390 6556 -241
rect 7292 -390 7313 -241
rect 7338 -390 7603 -371
rect 7626 -390 7647 -241
<< polysilicon >>
rect 4525 2737 4527 2739
rect 4535 2737 4537 2739
rect 4545 2737 4547 2739
rect 4555 2737 4557 2739
rect 4565 2737 4567 2739
rect 4575 2737 4577 2739
rect 4585 2737 4587 2739
rect 4595 2737 4597 2739
rect 4605 2737 4607 2739
rect 4615 2737 4617 2739
rect 4625 2737 4627 2739
rect 4635 2737 4637 2739
rect 4645 2737 4647 2739
rect 4450 2707 4452 2709
rect 4460 2707 4462 2709
rect 4470 2707 4472 2709
rect 4480 2707 4482 2709
rect 4425 2698 4427 2701
rect 4259 2658 4261 2660
rect 4297 2658 4299 2660
rect 4324 2658 4326 2660
rect 4347 2658 4349 2660
rect 4370 2658 4372 2660
rect 4259 2626 4261 2652
rect 4246 2624 4261 2626
rect 4259 2620 4261 2624
rect 4297 2620 4299 2652
rect 4324 2645 4326 2652
rect 4320 2643 4326 2645
rect 4259 2614 4261 2616
rect 4297 2610 4299 2616
rect 4246 2608 4299 2610
rect 4308 2610 4310 2623
rect 4324 2620 4326 2643
rect 4347 2620 4349 2652
rect 4370 2641 4372 2652
rect 4400 2651 4402 2653
rect 4361 2639 4372 2641
rect 4370 2620 4372 2639
rect 4655 2670 4657 2672
rect 4400 2630 4402 2637
rect 4397 2627 4402 2630
rect 4324 2614 4326 2616
rect 4347 2610 4349 2616
rect 4370 2614 4372 2616
rect 4400 2612 4402 2627
rect 4425 2630 4427 2637
rect 4422 2627 4427 2630
rect 4425 2615 4427 2627
rect 4450 2630 4452 2637
rect 4460 2630 4462 2637
rect 4470 2630 4472 2637
rect 4480 2630 4482 2637
rect 4447 2627 4482 2630
rect 4450 2615 4452 2627
rect 4460 2615 4462 2627
rect 4470 2615 4472 2627
rect 4480 2619 4482 2627
rect 4525 2630 4527 2637
rect 4535 2630 4537 2637
rect 4545 2630 4547 2637
rect 4555 2630 4557 2637
rect 4565 2630 4567 2637
rect 4575 2630 4577 2637
rect 4585 2630 4587 2637
rect 4595 2630 4597 2637
rect 4605 2630 4607 2637
rect 4615 2630 4617 2637
rect 4625 2630 4627 2637
rect 4635 2630 4637 2637
rect 4645 2630 4647 2637
rect 4655 2630 4657 2637
rect 4522 2627 4657 2630
rect 4480 2617 4502 2619
rect 4480 2615 4482 2617
rect 4490 2615 4492 2617
rect 4500 2615 4502 2617
rect 4525 2615 4527 2627
rect 4535 2615 4537 2627
rect 4545 2615 4547 2627
rect 4555 2615 4557 2627
rect 4565 2615 4567 2627
rect 4575 2615 4577 2627
rect 6584 2758 6586 2760
rect 6594 2758 6596 2760
rect 6604 2758 6606 2760
rect 6614 2758 6616 2760
rect 6624 2758 6626 2760
rect 6634 2758 6636 2760
rect 6644 2758 6646 2760
rect 6654 2758 6656 2760
rect 6664 2758 6666 2760
rect 6674 2758 6676 2760
rect 6684 2758 6686 2760
rect 6694 2758 6696 2760
rect 6704 2758 6706 2760
rect 6509 2728 6511 2730
rect 6519 2728 6521 2730
rect 6529 2728 6531 2730
rect 6539 2728 6541 2730
rect 6484 2719 6486 2722
rect 4308 2608 4349 2610
rect 4400 2604 4402 2606
rect 4500 2603 4502 2605
rect 4450 2593 4452 2595
rect 4460 2593 4462 2595
rect 4470 2593 4472 2595
rect 4480 2593 4482 2595
rect 4490 2593 4492 2595
rect 4425 2587 4427 2589
rect 6318 2679 6320 2681
rect 6356 2679 6358 2681
rect 6383 2679 6385 2681
rect 6406 2679 6408 2681
rect 6429 2679 6431 2681
rect 6318 2647 6320 2673
rect 6305 2645 6320 2647
rect 6318 2641 6320 2645
rect 6356 2641 6358 2673
rect 6383 2666 6385 2673
rect 6379 2664 6385 2666
rect 6318 2635 6320 2637
rect 6356 2631 6358 2637
rect 6305 2629 6358 2631
rect 6367 2631 6369 2644
rect 6383 2641 6385 2664
rect 6406 2641 6408 2673
rect 6429 2662 6431 2673
rect 6459 2672 6461 2674
rect 6420 2660 6431 2662
rect 6429 2641 6431 2660
rect 6714 2691 6716 2693
rect 6459 2651 6461 2658
rect 6456 2648 6461 2651
rect 6383 2635 6385 2637
rect 6406 2631 6408 2637
rect 6429 2635 6431 2637
rect 6459 2633 6461 2648
rect 6484 2651 6486 2658
rect 6481 2648 6486 2651
rect 6484 2636 6486 2648
rect 6509 2651 6511 2658
rect 6519 2651 6521 2658
rect 6529 2651 6531 2658
rect 6539 2651 6541 2658
rect 6506 2648 6541 2651
rect 6509 2636 6511 2648
rect 6519 2636 6521 2648
rect 6529 2636 6531 2648
rect 6539 2640 6541 2648
rect 6584 2651 6586 2658
rect 6594 2651 6596 2658
rect 6604 2651 6606 2658
rect 6614 2651 6616 2658
rect 6624 2651 6626 2658
rect 6634 2651 6636 2658
rect 6644 2651 6646 2658
rect 6654 2651 6656 2658
rect 6664 2651 6666 2658
rect 6674 2651 6676 2658
rect 6684 2651 6686 2658
rect 6694 2651 6696 2658
rect 6704 2651 6706 2658
rect 6714 2651 6716 2658
rect 6581 2648 6716 2651
rect 6539 2638 6561 2640
rect 6539 2636 6541 2638
rect 6549 2636 6551 2638
rect 6559 2636 6561 2638
rect 6584 2636 6586 2648
rect 6594 2636 6596 2648
rect 6604 2636 6606 2648
rect 6614 2636 6616 2648
rect 6624 2636 6626 2648
rect 6634 2636 6636 2648
rect 6367 2629 6408 2631
rect 6459 2625 6461 2627
rect 6559 2624 6561 2626
rect 6509 2614 6511 2616
rect 6519 2614 6521 2616
rect 6529 2614 6531 2616
rect 6539 2614 6541 2616
rect 6549 2614 6551 2616
rect 6484 2608 6486 2610
rect 4575 2558 4577 2560
rect 4525 2513 4527 2515
rect 4535 2513 4537 2515
rect 4545 2513 4547 2515
rect 4555 2513 4557 2515
rect 4565 2513 4567 2515
rect 6634 2579 6636 2581
rect 6584 2534 6586 2536
rect 6594 2534 6596 2536
rect 6604 2534 6606 2536
rect 6614 2534 6616 2536
rect 6624 2534 6626 2536
rect 4613 1155 4615 1157
rect 4623 1155 4625 1157
rect 4633 1155 4635 1157
rect 4643 1155 4645 1157
rect 4653 1155 4655 1157
rect 4603 1110 4605 1112
rect 6662 1127 6664 1129
rect 6672 1127 6674 1129
rect 6682 1127 6684 1129
rect 6692 1127 6694 1129
rect 6702 1127 6704 1129
rect 4753 1081 4755 1083
rect 4688 1075 4690 1077
rect 4698 1075 4700 1077
rect 4708 1075 4710 1077
rect 4718 1075 4720 1077
rect 4728 1075 4730 1077
rect 4678 1065 4680 1067
rect 4778 1064 4780 1066
rect 4831 1060 4872 1062
rect 4603 1043 4605 1055
rect 4613 1043 4615 1055
rect 4623 1043 4625 1055
rect 4633 1043 4635 1055
rect 4643 1043 4645 1055
rect 4653 1043 4655 1055
rect 4678 1053 4680 1055
rect 4688 1053 4690 1055
rect 4698 1053 4700 1055
rect 4678 1051 4700 1053
rect 4523 1040 4658 1043
rect 4523 1033 4525 1040
rect 4533 1033 4535 1040
rect 4543 1033 4545 1040
rect 4553 1033 4555 1040
rect 4563 1033 4565 1040
rect 4573 1033 4575 1040
rect 4583 1033 4585 1040
rect 4593 1033 4595 1040
rect 4603 1033 4605 1040
rect 4613 1033 4615 1040
rect 4623 1033 4625 1040
rect 4633 1033 4635 1040
rect 4643 1033 4645 1040
rect 4653 1033 4655 1040
rect 4698 1043 4700 1051
rect 4708 1043 4710 1055
rect 4718 1043 4720 1055
rect 4728 1043 4730 1055
rect 4698 1040 4733 1043
rect 4698 1033 4700 1040
rect 4708 1033 4710 1040
rect 4718 1033 4720 1040
rect 4728 1033 4730 1040
rect 4753 1043 4755 1055
rect 4753 1040 4758 1043
rect 4753 1033 4755 1040
rect 4778 1043 4780 1058
rect 4808 1054 4810 1056
rect 4831 1054 4833 1060
rect 4854 1054 4856 1056
rect 4778 1040 4783 1043
rect 4778 1033 4780 1040
rect 4523 998 4525 1000
rect 4808 1031 4810 1050
rect 4808 1029 4819 1031
rect 4778 1017 4780 1019
rect 4808 1018 4810 1029
rect 4831 1018 4833 1050
rect 4854 1027 4856 1050
rect 4870 1047 4872 1060
rect 4881 1060 4934 1062
rect 4881 1054 4883 1060
rect 4919 1054 4921 1056
rect 4854 1025 4860 1027
rect 4854 1018 4856 1025
rect 4881 1018 4883 1050
rect 4919 1046 4921 1050
rect 4919 1044 4934 1046
rect 4919 1018 4921 1044
rect 4808 1010 4810 1012
rect 4831 1010 4833 1012
rect 4854 1010 4856 1012
rect 4881 1010 4883 1012
rect 4919 1010 4921 1012
rect 6652 1082 6654 1084
rect 4753 969 4755 972
rect 4698 961 4700 963
rect 4708 961 4710 963
rect 4718 961 4720 963
rect 4728 961 4730 963
rect 4533 931 4535 933
rect 4543 931 4545 933
rect 4553 931 4555 933
rect 4563 931 4565 933
rect 4573 931 4575 933
rect 4583 931 4585 933
rect 4593 931 4595 933
rect 4603 931 4605 933
rect 4613 931 4615 933
rect 4623 931 4625 933
rect 4633 931 4635 933
rect 4643 931 4645 933
rect 4653 931 4655 933
rect 6802 1053 6804 1055
rect 6737 1047 6739 1049
rect 6747 1047 6749 1049
rect 6757 1047 6759 1049
rect 6767 1047 6769 1049
rect 6777 1047 6779 1049
rect 6727 1037 6729 1039
rect 6827 1036 6829 1038
rect 6880 1032 6921 1034
rect 6652 1015 6654 1027
rect 6662 1015 6664 1027
rect 6672 1015 6674 1027
rect 6682 1015 6684 1027
rect 6692 1015 6694 1027
rect 6702 1015 6704 1027
rect 6727 1025 6729 1027
rect 6737 1025 6739 1027
rect 6747 1025 6749 1027
rect 6727 1023 6749 1025
rect 6572 1012 6707 1015
rect 6572 1005 6574 1012
rect 6582 1005 6584 1012
rect 6592 1005 6594 1012
rect 6602 1005 6604 1012
rect 6612 1005 6614 1012
rect 6622 1005 6624 1012
rect 6632 1005 6634 1012
rect 6642 1005 6644 1012
rect 6652 1005 6654 1012
rect 6662 1005 6664 1012
rect 6672 1005 6674 1012
rect 6682 1005 6684 1012
rect 6692 1005 6694 1012
rect 6702 1005 6704 1012
rect 6747 1015 6749 1023
rect 6757 1015 6759 1027
rect 6767 1015 6769 1027
rect 6777 1015 6779 1027
rect 6747 1012 6782 1015
rect 6747 1005 6749 1012
rect 6757 1005 6759 1012
rect 6767 1005 6769 1012
rect 6777 1005 6779 1012
rect 6802 1015 6804 1027
rect 6802 1012 6807 1015
rect 6802 1005 6804 1012
rect 6827 1015 6829 1030
rect 6857 1026 6859 1028
rect 6880 1026 6882 1032
rect 6903 1026 6905 1028
rect 6827 1012 6832 1015
rect 6827 1005 6829 1012
rect 6572 970 6574 972
rect 6857 1003 6859 1022
rect 6857 1001 6868 1003
rect 6827 989 6829 991
rect 6857 990 6859 1001
rect 6880 990 6882 1022
rect 6903 999 6905 1022
rect 6919 1019 6921 1032
rect 6930 1032 6983 1034
rect 6930 1026 6932 1032
rect 6968 1026 6970 1028
rect 6903 997 6909 999
rect 6903 990 6905 997
rect 6930 990 6932 1022
rect 6968 1018 6970 1022
rect 6968 1016 6983 1018
rect 6968 990 6970 1016
rect 6857 982 6859 984
rect 6880 982 6882 984
rect 6903 982 6905 984
rect 6930 982 6932 984
rect 6968 982 6970 984
rect 6802 941 6804 944
rect 6747 933 6749 935
rect 6757 933 6759 935
rect 6767 933 6769 935
rect 6777 933 6779 935
rect 6582 903 6584 905
rect 6592 903 6594 905
rect 6602 903 6604 905
rect 6612 903 6614 905
rect 6622 903 6624 905
rect 6632 903 6634 905
rect 6642 903 6644 905
rect 6652 903 6654 905
rect 6662 903 6664 905
rect 6672 903 6674 905
rect 6682 903 6684 905
rect 6692 903 6694 905
rect 6702 903 6704 905
<< polycontact >>
rect 4241 2622 4246 2627
rect 4315 2642 4320 2647
rect 4306 2623 4311 2628
rect 4241 2606 4246 2611
rect 4356 2637 4361 2642
rect 4392 2626 4397 2631
rect 4417 2626 4422 2631
rect 4442 2626 4447 2631
rect 4517 2626 4522 2631
rect 6300 2643 6305 2648
rect 6374 2663 6379 2668
rect 6365 2644 6370 2649
rect 6300 2627 6305 2632
rect 6415 2658 6420 2663
rect 6451 2647 6456 2652
rect 6476 2647 6481 2652
rect 6501 2647 6506 2652
rect 6576 2647 6581 2652
rect 4658 1039 4663 1044
rect 4733 1039 4738 1044
rect 4758 1039 4763 1044
rect 4783 1039 4788 1044
rect 4819 1028 4824 1033
rect 4934 1059 4939 1064
rect 4869 1042 4874 1047
rect 4860 1023 4865 1028
rect 4934 1043 4939 1048
rect 6707 1011 6712 1016
rect 6782 1011 6787 1016
rect 6807 1011 6812 1016
rect 6832 1011 6837 1016
rect 6868 1000 6873 1005
rect 6983 1031 6988 1036
rect 6918 1014 6923 1019
rect 6909 995 6914 1000
rect 6983 1015 6988 1020
<< metal1 >>
rect 4984 4513 5050 4518
rect 4984 4511 5045 4513
rect 4984 4509 5043 4511
rect 4984 4507 5040 4509
rect 4985 4505 5038 4507
rect 7807 4506 7857 4509
rect 4987 4504 5038 4505
rect 7809 4504 7855 4506
rect 3781 4491 3873 4503
rect 4987 4502 5035 4504
rect 4989 4500 5033 4502
rect 4989 4499 5031 4500
rect 3788 4486 3866 4491
rect 3793 4479 3861 4486
rect 3800 4474 3854 4479
rect 3805 3682 3849 4474
rect 3907 3831 3930 3850
rect 4195 3831 4220 3850
rect 3927 3769 4196 3788
rect 4048 3682 4093 3769
rect 4992 3682 5031 4499
rect 6581 4498 6651 4503
rect 7812 4502 7852 4504
rect 7814 4499 7850 4502
rect 6586 4493 6646 4498
rect 7817 4497 7847 4499
rect 6591 4488 6641 4493
rect 6596 4483 6636 4488
rect 6601 4478 6631 4483
rect 5072 3831 5095 3850
rect 5360 3831 5385 3850
rect 5092 3769 5361 3788
rect 5213 3682 5258 3769
rect 6227 3831 6250 3850
rect 6515 3831 6540 3850
rect 6247 3769 6516 3788
rect 6368 3682 6413 3769
rect 6606 3682 6631 4478
rect 7420 3831 7443 3850
rect 7708 3831 7733 3850
rect 7440 3769 7709 3788
rect 7561 3682 7606 3769
rect 7819 3682 7845 4497
rect 3805 3680 4390 3682
rect 4745 3680 4760 3682
rect 3805 3608 4760 3680
rect 3805 3603 4423 3608
rect 3805 3600 4411 3603
rect 3805 3593 4390 3600
rect 4048 3525 4093 3593
rect 3929 3506 4196 3525
rect 3909 3436 3928 3457
rect 4203 3436 4222 3457
rect 4390 3375 4431 3444
rect 4738 3208 4760 3608
rect 4992 3593 5471 3682
rect 5213 3525 5258 3593
rect 5094 3506 5361 3525
rect 5074 3436 5093 3457
rect 5368 3436 5387 3457
rect 3238 2928 3865 2951
rect 3070 2820 3089 2845
rect 3070 2532 3089 2555
rect 3132 2718 3151 2821
rect 3238 2718 3327 2928
rect 3463 2828 3484 2847
rect 3395 2718 3414 2821
rect 3132 2673 3414 2718
rect 3132 2552 3151 2673
rect 2370 2473 2404 2479
rect 2370 2467 2409 2473
rect 2370 2462 2415 2467
rect 2370 2456 2421 2462
rect 3238 2456 3327 2673
rect 3395 2554 3414 2673
rect 3842 2646 3865 2928
rect 4745 2800 4760 3208
rect 4347 2779 4356 2785
rect 4362 2779 4365 2785
rect 4371 2779 4380 2785
rect 4347 2776 4353 2779
rect 4390 2771 4431 2790
rect 4437 2779 4446 2785
rect 4452 2779 4455 2785
rect 4461 2779 4464 2785
rect 4470 2779 4473 2785
rect 4479 2779 4482 2785
rect 4488 2779 4491 2785
rect 4497 2779 4500 2785
rect 4506 2779 4509 2785
rect 4515 2779 4518 2785
rect 4524 2779 4527 2785
rect 4533 2779 4536 2785
rect 4542 2779 4545 2785
rect 4551 2779 4554 2785
rect 4560 2779 4563 2785
rect 4569 2779 4572 2785
rect 4578 2779 4581 2785
rect 4587 2779 4590 2785
rect 4596 2779 4599 2785
rect 4605 2779 4608 2785
rect 4614 2779 4617 2785
rect 4623 2779 4626 2785
rect 4632 2779 4635 2785
rect 4641 2779 4644 2785
rect 4650 2779 4653 2785
rect 4659 2779 4662 2785
rect 4668 2779 4671 2785
rect 4677 2779 4680 2785
rect 4686 2779 4689 2785
rect 4695 2779 4704 2785
rect 4698 2776 4704 2779
rect 4347 2767 4353 2770
rect 4347 2758 4353 2761
rect 4347 2749 4353 2752
rect 4347 2741 4353 2743
rect 4347 2732 4353 2735
rect 4347 2723 4353 2726
rect 4347 2714 4353 2717
rect 4347 2705 4353 2708
rect 4347 2696 4353 2699
rect 4222 2690 4231 2696
rect 4237 2690 4240 2696
rect 4246 2690 4249 2696
rect 4255 2690 4258 2696
rect 4264 2690 4267 2696
rect 4273 2690 4276 2696
rect 4282 2690 4285 2696
rect 4291 2690 4294 2696
rect 4300 2690 4303 2696
rect 4309 2690 4312 2696
rect 4318 2690 4321 2696
rect 4327 2690 4330 2696
rect 4336 2690 4339 2696
rect 4345 2690 4353 2696
rect 4366 2765 4375 2771
rect 4381 2765 4384 2771
rect 4390 2765 4393 2771
rect 4399 2765 4402 2771
rect 4408 2765 4413 2771
rect 4419 2765 4422 2771
rect 4428 2765 4431 2771
rect 4437 2765 4440 2771
rect 4446 2765 4449 2771
rect 4455 2765 4460 2771
rect 4466 2765 4469 2771
rect 4475 2765 4478 2771
rect 4484 2765 4487 2771
rect 4493 2765 4496 2771
rect 4502 2765 4505 2771
rect 4511 2765 4514 2771
rect 4520 2765 4523 2771
rect 4529 2765 4532 2771
rect 4538 2765 4543 2771
rect 4549 2765 4552 2771
rect 4558 2765 4561 2771
rect 4567 2765 4570 2771
rect 4576 2765 4579 2771
rect 4585 2765 4590 2771
rect 4596 2765 4599 2771
rect 4605 2765 4608 2771
rect 4614 2765 4617 2771
rect 4623 2765 4626 2771
rect 4632 2765 4635 2771
rect 4641 2765 4644 2771
rect 4650 2765 4653 2771
rect 4659 2765 4662 2771
rect 4668 2765 4671 2771
rect 4677 2765 4686 2771
rect 4366 2762 4372 2765
rect 4366 2753 4372 2756
rect 4366 2744 4372 2747
rect 4366 2735 4372 2738
rect 4366 2727 4372 2729
rect 4366 2718 4372 2721
rect 4366 2709 4372 2712
rect 4366 2700 4372 2703
rect 4390 2755 4431 2765
rect 4680 2762 4686 2765
rect 4390 2743 4663 2755
rect 4390 2728 4513 2743
rect 4519 2737 4523 2743
rect 4539 2737 4543 2743
rect 4559 2737 4563 2743
rect 4579 2737 4583 2743
rect 4599 2737 4603 2743
rect 4619 2737 4623 2743
rect 4639 2737 4643 2743
rect 4390 2713 4509 2728
rect 4390 2700 4423 2713
rect 4366 2691 4372 2694
rect 4222 2688 4228 2690
rect 4366 2682 4372 2685
rect 4222 2679 4228 2682
rect 4222 2670 4228 2673
rect 4222 2661 4228 2664
rect 4222 2652 4228 2655
rect 3842 2641 4152 2646
rect 3842 2638 4154 2641
rect 3842 2633 4159 2638
rect 4222 2637 4228 2646
rect 4236 2676 4245 2682
rect 4251 2676 4254 2682
rect 4260 2676 4263 2682
rect 4269 2676 4272 2682
rect 4278 2676 4283 2682
rect 4289 2676 4292 2682
rect 4298 2676 4301 2682
rect 4307 2676 4310 2682
rect 4316 2676 4319 2682
rect 4325 2676 4330 2682
rect 4336 2676 4339 2682
rect 4345 2676 4348 2682
rect 4354 2676 4357 2682
rect 4363 2676 4372 2682
rect 4236 2670 4242 2676
rect 4394 2668 4398 2700
rect 4236 2661 4242 2664
rect 4236 2652 4242 2655
rect 4252 2663 4398 2668
rect 4252 2658 4257 2663
rect 4290 2658 4295 2663
rect 4317 2658 4322 2663
rect 4340 2658 4345 2663
rect 4363 2658 4368 2663
rect 4236 2637 4242 2646
rect 3842 2631 4162 2633
rect 3842 2628 4167 2631
rect 3842 2626 4169 2628
rect 3842 2623 4241 2626
rect 4263 2621 4268 2653
rect 4301 2621 4306 2653
rect 4315 2640 4320 2642
rect 4328 2642 4333 2653
rect 4351 2642 4356 2653
rect 4328 2637 4356 2642
rect 4317 2621 4322 2624
rect 4328 2621 4333 2637
rect 4374 2631 4379 2653
rect 4394 2651 4398 2663
rect 4419 2698 4423 2700
rect 4444 2707 4448 2713
rect 4464 2707 4468 2713
rect 4484 2712 4509 2713
rect 4484 2707 4488 2712
rect 4659 2670 4663 2743
rect 4680 2753 4686 2756
rect 4680 2744 4686 2747
rect 4680 2735 4686 2738
rect 4680 2726 4686 2729
rect 4680 2717 4686 2720
rect 4680 2708 4686 2711
rect 4680 2699 4686 2702
rect 4680 2690 4686 2693
rect 4680 2681 4686 2684
rect 4680 2672 4686 2675
rect 4680 2663 4686 2666
rect 4680 2654 4686 2657
rect 4680 2640 4686 2648
rect 4698 2767 4704 2770
rect 4698 2758 4704 2761
rect 4698 2749 4704 2752
rect 4698 2737 4704 2743
rect 4698 2728 4704 2731
rect 4698 2719 4704 2722
rect 4698 2710 4704 2713
rect 4698 2703 4704 2704
rect 4698 2694 4704 2697
rect 4698 2685 4704 2688
rect 4698 2676 4704 2679
rect 4698 2667 4704 2670
rect 4698 2658 4704 2661
rect 4698 2640 4704 2652
rect 4404 2631 4408 2637
rect 4429 2631 4433 2637
rect 4454 2631 4458 2637
rect 4474 2631 4478 2637
rect 4529 2631 4533 2637
rect 4549 2631 4553 2637
rect 4569 2631 4573 2637
rect 4589 2631 4593 2637
rect 4609 2631 4613 2637
rect 4629 2631 4633 2637
rect 4649 2631 4653 2637
rect 4745 2631 4757 2800
rect 4351 2621 4356 2624
rect 4374 2626 4392 2631
rect 4404 2626 4417 2631
rect 4429 2626 4442 2631
rect 4454 2626 4517 2631
rect 4529 2626 4757 2631
rect 5444 2640 5471 3593
rect 6125 3593 6631 3682
rect 7324 3593 7845 3682
rect 6125 2817 6148 3593
rect 6368 3525 6413 3593
rect 6249 3506 6516 3525
rect 6229 3436 6248 3457
rect 6523 3436 6542 3457
rect 6798 3377 6829 3441
rect 7561 3525 7606 3593
rect 7442 3506 7709 3525
rect 7422 3436 7441 3457
rect 7716 3436 7735 3457
rect 7737 2854 8204 2873
rect 6125 2805 6271 2817
rect 6260 2651 6271 2805
rect 6406 2800 6415 2806
rect 6421 2800 6424 2806
rect 6430 2800 6439 2806
rect 6406 2797 6412 2800
rect 6449 2792 6490 2811
rect 6496 2800 6505 2806
rect 6511 2800 6514 2806
rect 6520 2800 6523 2806
rect 6529 2800 6532 2806
rect 6538 2800 6541 2806
rect 6547 2800 6550 2806
rect 6556 2800 6559 2806
rect 6565 2800 6568 2806
rect 6574 2800 6577 2806
rect 6583 2800 6586 2806
rect 6592 2800 6595 2806
rect 6601 2800 6604 2806
rect 6610 2800 6613 2806
rect 6619 2800 6622 2806
rect 6628 2800 6631 2806
rect 6637 2800 6640 2806
rect 6646 2800 6649 2806
rect 6655 2800 6658 2806
rect 6664 2800 6667 2806
rect 6673 2800 6676 2806
rect 6682 2800 6685 2806
rect 6691 2800 6694 2806
rect 6700 2800 6703 2806
rect 6709 2800 6712 2806
rect 6718 2800 6721 2806
rect 6727 2800 6730 2806
rect 6736 2800 6739 2806
rect 6745 2800 6748 2806
rect 6754 2800 6763 2806
rect 6757 2797 6763 2800
rect 6406 2788 6412 2791
rect 6406 2779 6412 2782
rect 6406 2770 6412 2773
rect 6406 2762 6412 2764
rect 6406 2753 6412 2756
rect 6406 2744 6412 2747
rect 6406 2735 6412 2738
rect 6406 2726 6412 2729
rect 6406 2717 6412 2720
rect 6281 2711 6290 2717
rect 6296 2711 6299 2717
rect 6305 2711 6308 2717
rect 6314 2711 6317 2717
rect 6323 2711 6326 2717
rect 6332 2711 6335 2717
rect 6341 2711 6344 2717
rect 6350 2711 6353 2717
rect 6359 2711 6362 2717
rect 6368 2711 6371 2717
rect 6377 2711 6380 2717
rect 6386 2711 6389 2717
rect 6395 2711 6398 2717
rect 6404 2711 6412 2717
rect 6425 2786 6434 2792
rect 6440 2786 6443 2792
rect 6449 2786 6452 2792
rect 6458 2786 6461 2792
rect 6467 2786 6472 2792
rect 6478 2786 6481 2792
rect 6487 2786 6490 2792
rect 6496 2786 6499 2792
rect 6505 2786 6508 2792
rect 6514 2786 6519 2792
rect 6525 2786 6528 2792
rect 6534 2786 6537 2792
rect 6543 2786 6546 2792
rect 6552 2786 6555 2792
rect 6561 2786 6564 2792
rect 6570 2786 6573 2792
rect 6579 2786 6582 2792
rect 6588 2786 6591 2792
rect 6597 2786 6602 2792
rect 6608 2786 6611 2792
rect 6617 2786 6620 2792
rect 6626 2786 6629 2792
rect 6635 2786 6638 2792
rect 6644 2786 6649 2792
rect 6655 2786 6658 2792
rect 6664 2786 6667 2792
rect 6673 2786 6676 2792
rect 6682 2786 6685 2792
rect 6691 2786 6694 2792
rect 6700 2786 6703 2792
rect 6709 2786 6712 2792
rect 6718 2786 6721 2792
rect 6727 2786 6730 2792
rect 6736 2786 6745 2792
rect 6425 2783 6431 2786
rect 6425 2774 6431 2777
rect 6425 2765 6431 2768
rect 6425 2756 6431 2759
rect 6425 2748 6431 2750
rect 6425 2739 6431 2742
rect 6425 2730 6431 2733
rect 6425 2721 6431 2724
rect 6449 2776 6490 2786
rect 6739 2783 6745 2786
rect 6449 2764 6722 2776
rect 6449 2749 6572 2764
rect 6578 2758 6582 2764
rect 6598 2758 6602 2764
rect 6618 2758 6622 2764
rect 6638 2758 6642 2764
rect 6658 2758 6662 2764
rect 6678 2758 6682 2764
rect 6698 2758 6702 2764
rect 6449 2734 6568 2749
rect 6449 2721 6482 2734
rect 6425 2712 6431 2715
rect 6281 2709 6287 2711
rect 6425 2703 6431 2706
rect 6281 2700 6287 2703
rect 6281 2691 6287 2694
rect 6281 2682 6287 2685
rect 6281 2673 6287 2676
rect 6281 2658 6287 2667
rect 6295 2697 6304 2703
rect 6310 2697 6313 2703
rect 6319 2697 6322 2703
rect 6328 2697 6331 2703
rect 6337 2697 6342 2703
rect 6348 2697 6351 2703
rect 6357 2697 6360 2703
rect 6366 2697 6369 2703
rect 6375 2697 6378 2703
rect 6384 2697 6389 2703
rect 6395 2697 6398 2703
rect 6404 2697 6407 2703
rect 6413 2697 6416 2703
rect 6422 2697 6431 2703
rect 6295 2691 6301 2697
rect 6453 2689 6457 2721
rect 6295 2682 6301 2685
rect 6295 2673 6301 2676
rect 6311 2684 6457 2689
rect 6311 2679 6316 2684
rect 6349 2679 6354 2684
rect 6376 2679 6381 2684
rect 6399 2679 6404 2684
rect 6422 2679 6427 2684
rect 6295 2658 6301 2667
rect 6260 2650 6272 2651
rect 6260 2648 6274 2650
rect 6260 2647 6275 2648
rect 6260 2644 6300 2647
rect 6322 2642 6327 2674
rect 6360 2642 6365 2674
rect 6374 2661 6379 2663
rect 6387 2663 6392 2674
rect 6410 2663 6415 2674
rect 6387 2658 6415 2663
rect 5444 2639 6248 2640
rect 5444 2638 6251 2639
rect 5444 2637 6252 2638
rect 6376 2642 6381 2645
rect 6387 2642 6392 2658
rect 6433 2652 6438 2674
rect 6453 2672 6457 2684
rect 6478 2719 6482 2721
rect 6503 2728 6507 2734
rect 6523 2728 6527 2734
rect 6543 2733 6568 2734
rect 6543 2728 6547 2733
rect 6718 2691 6722 2764
rect 6739 2774 6745 2777
rect 6739 2765 6745 2768
rect 6739 2756 6745 2759
rect 6739 2747 6745 2750
rect 6739 2738 6745 2741
rect 6739 2729 6745 2732
rect 6739 2720 6745 2723
rect 6739 2711 6745 2714
rect 6739 2702 6745 2705
rect 6739 2693 6745 2696
rect 6739 2684 6745 2687
rect 6739 2675 6745 2678
rect 6739 2661 6745 2669
rect 6757 2788 6763 2791
rect 6757 2779 6763 2782
rect 6757 2770 6763 2773
rect 6757 2758 6763 2764
rect 6757 2749 6763 2752
rect 6757 2740 6763 2743
rect 6757 2731 6763 2734
rect 6757 2724 6763 2725
rect 6757 2715 6763 2718
rect 6757 2706 6763 2709
rect 6757 2697 6763 2700
rect 6757 2688 6763 2691
rect 6757 2679 6763 2682
rect 6757 2661 6763 2673
rect 6463 2652 6467 2658
rect 6488 2652 6492 2658
rect 6513 2652 6517 2658
rect 6533 2652 6537 2658
rect 6588 2652 6592 2658
rect 6608 2652 6612 2658
rect 6628 2652 6632 2658
rect 6648 2652 6652 2658
rect 6668 2652 6672 2658
rect 6688 2652 6692 2658
rect 6708 2652 6712 2658
rect 7737 2652 7747 2854
rect 7958 2776 7979 2795
rect 6410 2642 6415 2645
rect 6433 2647 6451 2652
rect 6463 2647 6476 2652
rect 6488 2647 6501 2652
rect 6513 2647 6576 2652
rect 6588 2647 7747 2652
rect 6433 2642 6438 2647
rect 5444 2635 6254 2637
rect 5444 2634 6255 2635
rect 5444 2633 6256 2634
rect 5444 2632 6258 2633
rect 6311 2632 6316 2637
rect 6349 2632 6354 2637
rect 6399 2632 6404 2637
rect 6422 2633 6427 2637
rect 6463 2633 6467 2647
rect 6488 2636 6492 2647
rect 6513 2636 6517 2647
rect 6533 2636 6537 2647
rect 6553 2636 6557 2647
rect 6588 2636 6592 2647
rect 6608 2636 6612 2647
rect 6628 2636 6632 2647
rect 6422 2632 6453 2633
rect 5444 2631 6259 2632
rect 5444 2628 6300 2631
rect 6311 2627 6453 2632
rect 4374 2621 4379 2626
rect 4252 2611 4257 2616
rect 4290 2611 4295 2616
rect 4340 2611 4345 2616
rect 4363 2612 4368 2616
rect 4404 2612 4408 2626
rect 4429 2615 4433 2626
rect 4454 2615 4458 2626
rect 4474 2615 4478 2626
rect 4494 2615 4498 2626
rect 4529 2615 4533 2626
rect 4549 2615 4553 2626
rect 4569 2615 4573 2626
rect 4363 2611 4394 2612
rect 3842 2607 4241 2610
rect 3842 2603 4166 2607
rect 4252 2606 4394 2611
rect 3842 2601 4162 2603
rect 3842 2597 4160 2601
rect 3842 2592 4156 2597
rect 3842 2587 4152 2592
rect 4222 2589 4228 2598
rect 4252 2589 4398 2606
rect 3463 2534 3484 2553
rect 2370 2410 3327 2456
rect 2370 2406 2419 2410
rect 2370 2399 2415 2406
rect 2370 2395 2409 2399
rect 2370 2389 2404 2395
rect 3842 2044 3865 2587
rect 4222 2581 4228 2583
rect 4375 2586 4398 2589
rect 4419 2586 4423 2589
rect 4444 2586 4448 2595
rect 4464 2586 4468 2595
rect 4484 2586 4488 2595
rect 4504 2586 4508 2605
rect 4222 2575 4231 2581
rect 4237 2575 4240 2581
rect 4246 2575 4249 2581
rect 4255 2575 4258 2581
rect 4264 2575 4267 2581
rect 4273 2575 4276 2581
rect 4282 2575 4285 2581
rect 4291 2575 4294 2581
rect 4300 2575 4303 2581
rect 4309 2575 4312 2581
rect 4318 2575 4321 2581
rect 4327 2575 4330 2581
rect 4336 2575 4339 2581
rect 4345 2575 4348 2581
rect 4354 2575 4355 2581
rect 4361 2575 4368 2581
rect 4362 2572 4368 2575
rect 4362 2563 4368 2566
rect 4375 2564 4508 2586
rect 4362 2556 4368 2557
rect 4362 2550 4371 2556
rect 4377 2550 4380 2556
rect 4386 2550 4389 2556
rect 4395 2550 4398 2556
rect 4404 2550 4407 2556
rect 4413 2550 4416 2556
rect 4422 2550 4425 2556
rect 4431 2550 4434 2556
rect 4440 2550 4443 2556
rect 4449 2550 4452 2556
rect 4458 2550 4461 2556
rect 4467 2550 4474 2556
rect 4468 2547 4474 2550
rect 4468 2538 4474 2541
rect 4468 2529 4474 2532
rect 4468 2520 4474 2523
rect 4468 2511 4474 2514
rect 4468 2502 4474 2505
rect 4468 2490 4474 2496
rect 4479 2506 4508 2564
rect 4519 2506 4523 2515
rect 4539 2506 4543 2515
rect 4559 2506 4563 2515
rect 4579 2506 4583 2560
rect 4479 2495 4583 2506
rect 4548 2490 4583 2495
rect 4600 2608 4609 2614
rect 4615 2608 4618 2614
rect 4624 2608 4627 2614
rect 4633 2608 4636 2614
rect 4642 2608 4645 2614
rect 4651 2608 4654 2614
rect 4660 2608 4663 2614
rect 4669 2608 4672 2614
rect 4678 2608 4681 2614
rect 4687 2608 4690 2614
rect 4696 2608 4704 2614
rect 6281 2610 6287 2619
rect 6311 2610 6457 2627
rect 4600 2605 4606 2608
rect 4600 2596 4606 2599
rect 6281 2602 6287 2604
rect 6434 2607 6457 2610
rect 6478 2607 6482 2610
rect 6503 2607 6507 2616
rect 6523 2607 6527 2616
rect 6543 2607 6547 2616
rect 6563 2607 6567 2626
rect 6281 2596 6290 2602
rect 6296 2596 6299 2602
rect 6305 2596 6308 2602
rect 6314 2596 6317 2602
rect 6323 2596 6326 2602
rect 6332 2596 6335 2602
rect 6341 2596 6344 2602
rect 6350 2596 6353 2602
rect 6359 2596 6362 2602
rect 6368 2596 6371 2602
rect 6377 2596 6380 2602
rect 6386 2596 6389 2602
rect 6395 2596 6398 2602
rect 6404 2596 6407 2602
rect 6413 2596 6414 2602
rect 6420 2596 6427 2602
rect 4600 2587 4606 2590
rect 4600 2578 4606 2581
rect 4600 2569 4606 2572
rect 6421 2593 6427 2596
rect 6421 2584 6427 2587
rect 6434 2585 6567 2607
rect 6421 2577 6427 2578
rect 6421 2571 6430 2577
rect 6436 2571 6439 2577
rect 6445 2571 6448 2577
rect 6454 2571 6457 2577
rect 6463 2571 6466 2577
rect 6472 2571 6475 2577
rect 6481 2571 6484 2577
rect 6490 2571 6493 2577
rect 6499 2571 6502 2577
rect 6508 2571 6511 2577
rect 6517 2571 6520 2577
rect 6526 2571 6533 2577
rect 4600 2560 4606 2563
rect 4600 2551 4606 2554
rect 4600 2542 4606 2545
rect 4600 2533 4606 2536
rect 4600 2524 4606 2527
rect 4600 2515 4606 2518
rect 4600 2506 4606 2509
rect 6527 2568 6533 2571
rect 6527 2559 6533 2562
rect 6527 2550 6533 2553
rect 6527 2541 6533 2544
rect 6527 2532 6533 2535
rect 6527 2523 6533 2526
rect 6527 2511 6533 2517
rect 6538 2527 6567 2585
rect 6578 2527 6582 2536
rect 6598 2527 6602 2536
rect 6618 2527 6622 2536
rect 6638 2527 6642 2581
rect 6538 2516 6642 2527
rect 6607 2511 6642 2516
rect 6659 2629 6668 2635
rect 6674 2629 6677 2635
rect 6683 2629 6686 2635
rect 6692 2629 6695 2635
rect 6701 2629 6704 2635
rect 6710 2629 6713 2635
rect 6719 2629 6722 2635
rect 6728 2629 6731 2635
rect 6737 2629 6740 2635
rect 6746 2629 6749 2635
rect 6755 2629 6763 2635
rect 6659 2626 6665 2629
rect 6659 2617 6665 2620
rect 6659 2608 6665 2611
rect 6659 2599 6665 2602
rect 6659 2590 6665 2593
rect 6659 2581 6665 2584
rect 6659 2572 6665 2575
rect 6659 2563 6665 2566
rect 6659 2554 6665 2557
rect 6659 2545 6665 2548
rect 6659 2536 6665 2539
rect 6659 2527 6665 2530
rect 6659 2518 6665 2521
rect 6527 2505 6536 2511
rect 6542 2505 6545 2511
rect 6551 2505 6554 2511
rect 6560 2505 6563 2511
rect 6569 2505 6572 2511
rect 6578 2505 6581 2511
rect 6587 2505 6590 2511
rect 6596 2505 6599 2511
rect 6605 2505 6608 2511
rect 6614 2505 6617 2511
rect 6623 2505 6626 2511
rect 6632 2505 6635 2511
rect 6641 2505 6644 2511
rect 6650 2505 6653 2511
rect 6659 2505 6665 2512
rect 4600 2497 4606 2500
rect 4468 2484 4477 2490
rect 4483 2484 4486 2490
rect 4492 2484 4495 2490
rect 4501 2484 4504 2490
rect 4510 2484 4513 2490
rect 4519 2484 4522 2490
rect 4528 2484 4531 2490
rect 4537 2484 4540 2490
rect 4546 2484 4549 2490
rect 4555 2484 4558 2490
rect 4564 2484 4567 2490
rect 4573 2484 4576 2490
rect 4582 2484 4585 2490
rect 4591 2484 4594 2490
rect 4600 2484 4606 2491
rect 6607 2496 6642 2505
rect 8028 2656 8047 2775
rect 8115 2656 8204 2854
rect 8291 2656 8310 2777
rect 8028 2611 8310 2656
rect 8028 2508 8047 2611
rect 4548 2475 4583 2484
rect 7958 2482 7979 2501
rect 8115 2409 8204 2611
rect 8291 2508 8310 2611
rect 8353 2774 8372 2797
rect 8353 2484 8372 2509
rect 9063 2429 9067 2433
rect 9056 2423 9067 2429
rect 9052 2419 9067 2423
rect 9045 2413 9067 2419
rect 9041 2409 9067 2413
rect 8115 2383 9067 2409
rect 9041 2379 9067 2383
rect 9045 2373 9067 2379
rect 9052 2369 9067 2373
rect 9056 2363 9067 2369
rect 9063 2359 9067 2363
rect 9070 2067 9073 2068
rect 9068 2065 9073 2067
rect 9067 2064 9073 2065
rect 9065 2062 9073 2064
rect 9064 2061 9073 2062
rect 9062 2059 9073 2061
rect 9061 2058 9073 2059
rect 9059 2056 9073 2058
rect 9058 2055 9073 2056
rect 9056 2053 9073 2055
rect 3237 2021 3865 2044
rect 8115 2030 9073 2053
rect 3069 1910 3088 1935
rect 3069 1622 3088 1645
rect 3131 1808 3150 1911
rect 3237 1808 3326 2021
rect 3462 1918 3483 1937
rect 7958 1930 7979 1949
rect 3394 1808 3413 1911
rect 3131 1763 3413 1808
rect 3131 1642 3150 1763
rect 2368 1597 2402 1603
rect 3237 1603 3326 1763
rect 3394 1644 3413 1763
rect 8028 1810 8047 1929
rect 8115 1810 8204 2030
rect 9056 2028 9073 2030
rect 9058 2027 9073 2028
rect 9059 2025 9073 2027
rect 9061 2024 9073 2025
rect 9062 2022 9073 2024
rect 9064 2021 9073 2022
rect 9065 2019 9073 2021
rect 9067 2018 9073 2019
rect 9068 2016 9073 2018
rect 9070 2015 9073 2016
rect 8291 1810 8310 1931
rect 8028 1765 8310 1810
rect 8028 1662 8047 1765
rect 3462 1624 3483 1643
rect 2368 1591 2407 1597
rect 2368 1586 2413 1591
rect 2368 1580 2419 1586
rect 3236 1580 3326 1603
rect 7958 1636 7979 1655
rect 2368 1542 3326 1580
rect 8115 1552 8204 1765
rect 8291 1662 8310 1765
rect 8353 1928 8372 1951
rect 8353 1638 8372 1663
rect 2368 1534 3325 1542
rect 2368 1530 2417 1534
rect 2368 1523 2413 1530
rect 2368 1519 2407 1523
rect 2368 1513 2402 1519
rect 8140 1373 8175 1552
rect 8139 1294 8175 1373
rect 7831 1266 8175 1294
rect 4597 1186 4632 1195
rect 4574 1179 4580 1186
rect 4586 1180 4589 1186
rect 4595 1180 4598 1186
rect 4604 1180 4607 1186
rect 4613 1180 4616 1186
rect 4622 1180 4625 1186
rect 4631 1180 4634 1186
rect 4640 1180 4643 1186
rect 4649 1180 4652 1186
rect 4658 1180 4661 1186
rect 4667 1180 4670 1186
rect 4676 1180 4679 1186
rect 4685 1180 4688 1186
rect 4694 1180 4697 1186
rect 4703 1180 4712 1186
rect 4574 1170 4580 1173
rect 4574 1161 4580 1164
rect 4574 1152 4580 1155
rect 4574 1143 4580 1146
rect 4574 1134 4580 1137
rect 4574 1125 4580 1128
rect 4574 1116 4580 1119
rect 4574 1107 4580 1110
rect 4574 1098 4580 1101
rect 2374 1094 2377 1096
rect 2374 1091 2379 1094
rect 2374 1089 2381 1091
rect 4574 1089 4580 1092
rect 2374 1086 2384 1089
rect 2374 1084 2386 1086
rect 2374 1059 3326 1084
rect 4574 1080 4580 1083
rect 4574 1071 4580 1074
rect 4574 1062 4580 1065
rect 2374 1057 2386 1059
rect 2374 1054 2384 1057
rect 2374 1052 2381 1054
rect 2374 1049 2379 1052
rect 2374 1047 2377 1049
rect 3069 970 3088 995
rect 3069 682 3088 705
rect 3131 868 3150 971
rect 3237 868 3326 1059
rect 4476 1056 4484 1062
rect 4490 1056 4493 1062
rect 4499 1056 4502 1062
rect 4508 1056 4511 1062
rect 4517 1056 4520 1062
rect 4526 1056 4529 1062
rect 4535 1056 4538 1062
rect 4544 1056 4547 1062
rect 4553 1056 4556 1062
rect 4562 1056 4565 1062
rect 4571 1056 4580 1062
rect 4597 1175 4632 1180
rect 4597 1164 4701 1175
rect 4597 1110 4601 1164
rect 4617 1155 4621 1164
rect 4637 1155 4641 1164
rect 4657 1155 4661 1164
rect 4672 1106 4701 1164
rect 4706 1174 4712 1180
rect 4706 1165 4712 1168
rect 4706 1156 4712 1159
rect 6646 1158 6681 1167
rect 4706 1147 4712 1150
rect 4706 1138 4712 1141
rect 4706 1129 4712 1132
rect 4706 1120 4712 1123
rect 6623 1151 6629 1158
rect 6635 1152 6638 1158
rect 6644 1152 6647 1158
rect 6653 1152 6656 1158
rect 6662 1152 6665 1158
rect 6671 1152 6674 1158
rect 6680 1152 6683 1158
rect 6689 1152 6692 1158
rect 6698 1152 6701 1158
rect 6707 1152 6710 1158
rect 6716 1152 6719 1158
rect 6725 1152 6728 1158
rect 6734 1152 6737 1158
rect 6743 1152 6746 1158
rect 6752 1152 6761 1158
rect 6623 1142 6629 1145
rect 6623 1133 6629 1136
rect 6623 1124 6629 1127
rect 4706 1114 4713 1120
rect 4719 1114 4722 1120
rect 4728 1114 4731 1120
rect 4737 1114 4740 1120
rect 4746 1114 4749 1120
rect 4755 1114 4758 1120
rect 4764 1114 4767 1120
rect 4773 1114 4776 1120
rect 4782 1114 4785 1120
rect 4791 1114 4794 1120
rect 4800 1114 4803 1120
rect 4809 1114 4818 1120
rect 4812 1113 4818 1114
rect 4672 1084 4805 1106
rect 4812 1104 4818 1107
rect 4812 1095 4818 1098
rect 6623 1115 6629 1118
rect 6623 1106 6629 1109
rect 6623 1097 6629 1100
rect 4812 1089 4819 1095
rect 4825 1089 4826 1095
rect 4832 1089 4835 1095
rect 4841 1089 4844 1095
rect 4850 1089 4853 1095
rect 4859 1089 4862 1095
rect 4868 1089 4871 1095
rect 4877 1089 4880 1095
rect 4886 1089 4889 1095
rect 4895 1089 4898 1095
rect 4904 1089 4907 1095
rect 4913 1089 4916 1095
rect 4922 1089 4925 1095
rect 4931 1089 4934 1095
rect 4940 1089 4943 1095
rect 4949 1089 4958 1095
rect 4672 1065 4676 1084
rect 4692 1075 4696 1084
rect 4712 1075 4716 1084
rect 4732 1075 4736 1084
rect 4757 1081 4761 1084
rect 4782 1081 4805 1084
rect 4952 1087 4958 1089
rect 4782 1064 4928 1081
rect 4952 1072 4958 1081
rect 6623 1088 6629 1091
rect 6623 1079 6629 1082
rect 6623 1070 6629 1073
rect 4786 1059 4928 1064
rect 4939 1060 5049 1063
rect 4786 1058 4817 1059
rect 3717 1046 4464 1047
rect 3717 1045 4467 1046
rect 3717 1044 4470 1045
rect 4607 1044 4611 1055
rect 4627 1044 4631 1055
rect 4647 1044 4651 1055
rect 4682 1044 4686 1055
rect 4702 1044 4706 1055
rect 4722 1044 4726 1055
rect 4747 1044 4751 1055
rect 4772 1044 4776 1058
rect 4812 1054 4817 1058
rect 4835 1054 4840 1059
rect 4885 1054 4890 1059
rect 4923 1054 4928 1059
rect 4801 1044 4806 1049
rect 3717 1039 4651 1044
rect 4663 1039 4726 1044
rect 4738 1039 4751 1044
rect 4763 1039 4776 1044
rect 4788 1039 4806 1044
rect 4824 1046 4829 1049
rect 3717 1038 4470 1039
rect 3717 1037 4467 1038
rect 3717 1036 4464 1037
rect 3717 1034 4462 1036
rect 3717 1033 4460 1034
rect 4527 1033 4531 1039
rect 4547 1033 4551 1039
rect 4567 1033 4571 1039
rect 4587 1033 4591 1039
rect 4607 1033 4611 1039
rect 4627 1033 4631 1039
rect 4647 1033 4651 1039
rect 4702 1033 4706 1039
rect 4722 1033 4726 1039
rect 4747 1033 4751 1039
rect 4772 1033 4776 1039
rect 3717 1032 4457 1033
rect 3717 1031 4455 1032
rect 3717 1030 4452 1031
rect 3717 1029 4450 1030
rect 3717 1028 4446 1029
rect 3462 978 3483 997
rect 3394 868 3413 971
rect 3131 823 3413 868
rect 3131 702 3150 823
rect 3237 625 3326 823
rect 3394 704 3413 823
rect 3462 684 3483 703
rect 3717 625 3736 1028
rect 4476 1018 4482 1030
rect 4476 1009 4482 1012
rect 4476 1000 4482 1003
rect 4476 991 4482 994
rect 4476 982 4482 985
rect 4476 973 4482 976
rect 4476 966 4482 967
rect 4476 957 4482 960
rect 4476 948 4482 951
rect 4476 939 4482 942
rect 4476 927 4482 933
rect 4476 918 4482 921
rect 4476 909 4482 912
rect 4476 900 4482 903
rect 4494 1022 4500 1030
rect 4494 1013 4500 1016
rect 4494 1004 4500 1007
rect 4494 995 4500 998
rect 4494 986 4500 989
rect 4494 977 4500 980
rect 4494 968 4500 971
rect 4494 959 4500 962
rect 4494 950 4500 953
rect 4494 941 4500 944
rect 4494 932 4500 935
rect 4494 923 4500 926
rect 4494 914 4500 917
rect 4517 927 4521 1000
rect 4692 958 4696 963
rect 4671 957 4696 958
rect 4712 957 4716 963
rect 4732 957 4736 963
rect 4757 970 4761 972
rect 4782 1007 4786 1019
rect 4801 1017 4806 1039
rect 4847 1033 4852 1049
rect 4858 1046 4863 1049
rect 4824 1028 4852 1033
rect 4824 1017 4829 1028
rect 4847 1017 4852 1028
rect 4860 1028 4865 1030
rect 4874 1017 4879 1049
rect 4912 1017 4917 1049
rect 4968 1047 4999 1048
rect 4939 1044 4999 1047
rect 4938 1024 4944 1033
rect 4812 1007 4817 1012
rect 4835 1007 4840 1012
rect 4858 1007 4863 1012
rect 4885 1007 4890 1012
rect 4923 1007 4928 1012
rect 4782 1002 4928 1007
rect 4938 1015 4944 1018
rect 4938 1006 4944 1009
rect 4782 970 4786 1002
rect 4938 994 4944 1000
rect 4808 988 4817 994
rect 4823 988 4826 994
rect 4832 988 4835 994
rect 4841 988 4844 994
rect 4850 988 4855 994
rect 4861 988 4864 994
rect 4870 988 4873 994
rect 4879 988 4882 994
rect 4888 988 4891 994
rect 4897 988 4902 994
rect 4908 988 4911 994
rect 4917 988 4920 994
rect 4926 988 4929 994
rect 4935 988 4944 994
rect 4952 1024 4958 1033
rect 4952 1015 4958 1018
rect 4952 1006 4958 1009
rect 4952 997 4958 1000
rect 4952 988 4958 991
rect 4808 985 4814 988
rect 4952 980 4958 982
rect 4808 976 4814 979
rect 4757 957 4790 970
rect 4671 942 4790 957
rect 4537 927 4541 933
rect 4557 927 4561 933
rect 4577 927 4581 933
rect 4597 927 4601 933
rect 4617 927 4621 933
rect 4637 927 4641 933
rect 4657 927 4661 933
rect 4667 927 4790 942
rect 4517 915 4790 927
rect 4494 905 4500 908
rect 4749 905 4790 915
rect 4808 967 4814 970
rect 4808 958 4814 961
rect 4808 949 4814 952
rect 4808 941 4814 943
rect 4808 932 4814 935
rect 4808 923 4814 926
rect 4808 914 4814 917
rect 4808 905 4814 908
rect 4494 899 4503 905
rect 4509 899 4512 905
rect 4518 899 4521 905
rect 4527 899 4530 905
rect 4536 899 4539 905
rect 4545 899 4548 905
rect 4554 899 4557 905
rect 4563 899 4566 905
rect 4572 899 4575 905
rect 4581 899 4584 905
rect 4590 899 4595 905
rect 4601 899 4604 905
rect 4610 899 4613 905
rect 4619 899 4622 905
rect 4628 899 4631 905
rect 4637 899 4642 905
rect 4648 899 4651 905
rect 4657 899 4660 905
rect 4666 899 4669 905
rect 4675 899 4678 905
rect 4684 899 4687 905
rect 4693 899 4696 905
rect 4702 899 4705 905
rect 4711 899 4714 905
rect 4720 899 4725 905
rect 4731 899 4734 905
rect 4740 899 4743 905
rect 4749 899 4752 905
rect 4758 899 4761 905
rect 4767 899 4772 905
rect 4778 899 4781 905
rect 4787 899 4790 905
rect 4796 899 4799 905
rect 4805 899 4808 905
rect 4827 974 4835 980
rect 4841 974 4844 980
rect 4850 974 4853 980
rect 4859 974 4862 980
rect 4868 974 4871 980
rect 4877 974 4880 980
rect 4886 974 4889 980
rect 4895 974 4898 980
rect 4904 974 4907 980
rect 4913 974 4916 980
rect 4922 974 4925 980
rect 4931 974 4934 980
rect 4940 974 4943 980
rect 4949 974 4958 980
rect 4827 971 4833 974
rect 4827 962 4833 965
rect 4827 953 4833 956
rect 4827 944 4833 947
rect 4827 935 4833 938
rect 4827 927 4833 929
rect 4827 918 4833 921
rect 4827 909 4833 912
rect 4827 900 4833 903
rect 4476 891 4482 894
rect 4476 885 4485 891
rect 4491 885 4494 891
rect 4500 885 4503 891
rect 4509 885 4512 891
rect 4518 885 4521 891
rect 4527 885 4530 891
rect 4536 885 4539 891
rect 4545 885 4548 891
rect 4554 885 4557 891
rect 4563 885 4566 891
rect 4572 885 4575 891
rect 4581 885 4584 891
rect 4590 885 4593 891
rect 4599 885 4602 891
rect 4608 885 4611 891
rect 4617 885 4620 891
rect 4626 885 4629 891
rect 4635 885 4638 891
rect 4644 885 4647 891
rect 4653 885 4656 891
rect 4662 885 4665 891
rect 4671 885 4674 891
rect 4680 885 4683 891
rect 4689 885 4692 891
rect 4698 885 4701 891
rect 4707 885 4710 891
rect 4716 885 4719 891
rect 4725 885 4728 891
rect 4734 885 4743 891
rect 4749 880 4790 899
rect 4827 891 4833 894
rect 4800 885 4809 891
rect 4815 885 4818 891
rect 4824 885 4833 891
rect 4980 848 4999 1044
rect 3237 606 3736 625
rect 3831 823 4999 848
rect 3831 -134 3855 823
rect 5030 803 5049 1060
rect 6623 1061 6629 1064
rect 6623 1052 6629 1055
rect 6623 1043 6629 1046
rect 6623 1034 6629 1037
rect 6525 1028 6533 1034
rect 6539 1028 6542 1034
rect 6548 1028 6551 1034
rect 6557 1028 6560 1034
rect 6566 1028 6569 1034
rect 6575 1028 6578 1034
rect 6584 1028 6587 1034
rect 6593 1028 6596 1034
rect 6602 1028 6605 1034
rect 6611 1028 6614 1034
rect 6620 1028 6629 1034
rect 6646 1147 6681 1152
rect 6646 1136 6750 1147
rect 6646 1082 6650 1136
rect 6666 1127 6670 1136
rect 6686 1127 6690 1136
rect 6706 1127 6710 1136
rect 6721 1078 6750 1136
rect 6755 1146 6761 1152
rect 6755 1137 6761 1140
rect 6755 1128 6761 1131
rect 6755 1119 6761 1122
rect 6755 1110 6761 1113
rect 6755 1101 6761 1104
rect 6755 1092 6761 1095
rect 6755 1086 6762 1092
rect 6768 1086 6771 1092
rect 6777 1086 6780 1092
rect 6786 1086 6789 1092
rect 6795 1086 6798 1092
rect 6804 1086 6807 1092
rect 6813 1086 6816 1092
rect 6822 1086 6825 1092
rect 6831 1086 6834 1092
rect 6840 1086 6843 1092
rect 6849 1086 6852 1092
rect 6858 1086 6867 1092
rect 6861 1085 6867 1086
rect 6721 1056 6854 1078
rect 6861 1076 6867 1079
rect 6861 1067 6867 1070
rect 6861 1061 6868 1067
rect 6874 1061 6875 1067
rect 6881 1061 6884 1067
rect 6890 1061 6893 1067
rect 6899 1061 6902 1067
rect 6908 1061 6911 1067
rect 6917 1061 6920 1067
rect 6926 1061 6929 1067
rect 6935 1061 6938 1067
rect 6944 1061 6947 1067
rect 6953 1061 6956 1067
rect 6962 1061 6965 1067
rect 6971 1061 6974 1067
rect 6980 1061 6983 1067
rect 6989 1061 6992 1067
rect 6998 1061 7007 1067
rect 6721 1037 6725 1056
rect 6741 1047 6745 1056
rect 6761 1047 6765 1056
rect 6781 1047 6785 1056
rect 6806 1053 6810 1056
rect 6831 1053 6854 1056
rect 7001 1059 7007 1061
rect 6831 1036 6977 1053
rect 7001 1044 7007 1053
rect 7831 1043 7866 1266
rect 7081 1042 7866 1043
rect 7078 1041 7866 1042
rect 7075 1039 7866 1041
rect 7020 1038 7866 1039
rect 6835 1031 6977 1036
rect 7017 1035 7866 1038
rect 6988 1032 7866 1035
rect 6835 1030 6866 1031
rect 6656 1016 6660 1027
rect 6676 1016 6680 1027
rect 6696 1016 6700 1027
rect 6731 1016 6735 1027
rect 6751 1016 6755 1027
rect 6771 1016 6775 1027
rect 6796 1016 6800 1027
rect 6821 1016 6825 1030
rect 6861 1026 6866 1030
rect 6884 1026 6889 1031
rect 6934 1026 6939 1031
rect 6972 1026 6977 1031
rect 6850 1016 6855 1021
rect 4985 787 5049 803
rect 6130 1011 6700 1016
rect 6712 1011 6775 1016
rect 6787 1011 6800 1016
rect 6812 1011 6825 1016
rect 6837 1011 6855 1016
rect 6873 1018 6878 1021
rect 6130 1008 6502 1011
rect 6130 1006 6432 1008
rect 6130 1002 6365 1006
rect 6576 1005 6580 1011
rect 6596 1005 6600 1011
rect 6616 1005 6620 1011
rect 6636 1005 6640 1011
rect 6656 1005 6660 1011
rect 6676 1005 6680 1011
rect 6696 1005 6700 1011
rect 6751 1005 6755 1011
rect 6771 1005 6775 1011
rect 6796 1005 6800 1011
rect 6821 1005 6825 1011
rect 3915 2 3934 23
rect 4209 2 4228 23
rect 3941 -66 4208 -47
rect 4044 -134 4089 -66
rect 4749 10 4790 108
rect 4985 -133 5009 787
rect 5069 3 5088 24
rect 5363 3 5382 24
rect 5095 -65 5362 -46
rect 5198 -133 5243 -65
rect 6130 -133 6153 1002
rect 6525 990 6531 1002
rect 6525 981 6531 984
rect 6525 972 6531 975
rect 6525 963 6531 966
rect 6525 954 6531 957
rect 6525 945 6531 948
rect 6525 938 6531 939
rect 6525 929 6531 932
rect 6525 920 6531 923
rect 6525 911 6531 914
rect 6525 899 6531 905
rect 6525 890 6531 893
rect 6525 881 6531 884
rect 6525 872 6531 875
rect 6543 994 6549 1002
rect 6543 985 6549 988
rect 6543 976 6549 979
rect 6543 967 6549 970
rect 6543 958 6549 961
rect 6543 949 6549 952
rect 6543 940 6549 943
rect 6543 931 6549 934
rect 6543 922 6549 925
rect 6543 913 6549 916
rect 6543 904 6549 907
rect 6543 895 6549 898
rect 6543 886 6549 889
rect 6566 899 6570 972
rect 6741 930 6745 935
rect 6720 929 6745 930
rect 6761 929 6765 935
rect 6781 929 6785 935
rect 6806 942 6810 944
rect 6831 979 6835 991
rect 6850 989 6855 1011
rect 6896 1005 6901 1021
rect 6907 1018 6912 1021
rect 6873 1000 6901 1005
rect 6873 989 6878 1000
rect 6896 989 6901 1000
rect 6909 1000 6914 1002
rect 6923 989 6928 1021
rect 6961 989 6966 1021
rect 6988 1016 8203 1019
rect 7097 1015 8203 1016
rect 7098 1014 8203 1015
rect 7099 1013 8203 1014
rect 7100 1012 8203 1013
rect 7371 1010 8203 1012
rect 7373 1009 8203 1010
rect 7376 1008 8203 1009
rect 6987 996 6993 1005
rect 6861 979 6866 984
rect 6884 979 6889 984
rect 6907 979 6912 984
rect 6934 979 6939 984
rect 6972 979 6977 984
rect 6831 974 6977 979
rect 6987 987 6993 990
rect 6987 978 6993 981
rect 6831 942 6835 974
rect 6987 966 6993 972
rect 6857 960 6866 966
rect 6872 960 6875 966
rect 6881 960 6884 966
rect 6890 960 6893 966
rect 6899 960 6904 966
rect 6910 960 6913 966
rect 6919 960 6922 966
rect 6928 960 6931 966
rect 6937 960 6940 966
rect 6946 960 6951 966
rect 6957 960 6960 966
rect 6966 960 6969 966
rect 6975 960 6978 966
rect 6984 960 6993 966
rect 7001 996 7007 1005
rect 7001 987 7007 990
rect 7001 978 7007 981
rect 7001 969 7007 972
rect 7001 960 7007 963
rect 6857 957 6863 960
rect 7001 952 7007 954
rect 6857 948 6863 951
rect 6806 929 6839 942
rect 6720 914 6839 929
rect 6586 899 6590 905
rect 6606 899 6610 905
rect 6626 899 6630 905
rect 6646 899 6650 905
rect 6666 899 6670 905
rect 6686 899 6690 905
rect 6706 899 6710 905
rect 6716 899 6839 914
rect 6566 887 6839 899
rect 6543 877 6549 880
rect 6798 877 6839 887
rect 6857 939 6863 942
rect 6857 930 6863 933
rect 6857 921 6863 924
rect 6857 913 6863 915
rect 6857 904 6863 907
rect 6857 895 6863 898
rect 6857 886 6863 889
rect 6857 877 6863 880
rect 6543 871 6552 877
rect 6558 871 6561 877
rect 6567 871 6570 877
rect 6576 871 6579 877
rect 6585 871 6588 877
rect 6594 871 6597 877
rect 6603 871 6606 877
rect 6612 871 6615 877
rect 6621 871 6624 877
rect 6630 871 6633 877
rect 6639 871 6644 877
rect 6650 871 6653 877
rect 6659 871 6662 877
rect 6668 871 6671 877
rect 6677 871 6680 877
rect 6686 871 6691 877
rect 6697 871 6700 877
rect 6706 871 6709 877
rect 6715 871 6718 877
rect 6724 871 6727 877
rect 6733 871 6736 877
rect 6742 871 6745 877
rect 6751 871 6754 877
rect 6760 871 6763 877
rect 6769 871 6774 877
rect 6780 871 6783 877
rect 6789 871 6792 877
rect 6798 871 6801 877
rect 6807 871 6810 877
rect 6816 871 6821 877
rect 6827 871 6830 877
rect 6836 871 6839 877
rect 6845 871 6848 877
rect 6854 871 6863 877
rect 6876 946 6884 952
rect 6890 946 6893 952
rect 6899 946 6902 952
rect 6908 946 6911 952
rect 6917 946 6920 952
rect 6926 946 6929 952
rect 6935 946 6938 952
rect 6944 946 6947 952
rect 6953 946 6956 952
rect 6962 946 6965 952
rect 6971 946 6974 952
rect 6980 946 6983 952
rect 6989 946 6992 952
rect 6998 946 7007 952
rect 6876 943 6882 946
rect 6876 934 6882 937
rect 6876 925 6882 928
rect 6876 916 6882 919
rect 6876 907 6882 910
rect 7957 926 7978 945
rect 6876 899 6882 901
rect 6876 890 6882 893
rect 6876 881 6882 884
rect 6876 872 6882 875
rect 6525 863 6531 866
rect 6525 857 6534 863
rect 6540 857 6543 863
rect 6549 857 6552 863
rect 6558 857 6561 863
rect 6567 857 6570 863
rect 6576 857 6579 863
rect 6585 857 6588 863
rect 6594 857 6597 863
rect 6603 857 6606 863
rect 6612 857 6615 863
rect 6621 857 6624 863
rect 6630 857 6633 863
rect 6639 857 6642 863
rect 6648 857 6651 863
rect 6657 857 6660 863
rect 6666 857 6669 863
rect 6675 857 6678 863
rect 6684 857 6687 863
rect 6693 857 6696 863
rect 6702 857 6705 863
rect 6711 857 6714 863
rect 6720 857 6723 863
rect 6729 857 6732 863
rect 6738 857 6741 863
rect 6747 857 6750 863
rect 6756 857 6759 863
rect 6765 857 6768 863
rect 6774 857 6777 863
rect 6783 857 6792 863
rect 6798 852 6839 871
rect 6876 863 6882 866
rect 6855 857 6858 863
rect 6864 857 6867 863
rect 6873 857 6882 863
rect 8027 806 8046 925
rect 8114 806 8203 1008
rect 8290 806 8309 927
rect 8027 761 8309 806
rect 8027 658 8046 761
rect 7957 632 7978 651
rect 8114 562 8203 761
rect 8290 658 8309 761
rect 8352 924 8371 947
rect 8352 634 8371 659
rect 9068 569 9071 572
rect 9066 567 9071 569
rect 9063 564 9071 567
rect 9061 563 9071 564
rect 9059 562 9071 563
rect 8114 541 9071 562
rect 9063 540 9071 541
rect 9066 538 9071 540
rect 9068 535 9071 538
rect 6220 3 6239 24
rect 6514 3 6533 24
rect 6246 -65 6513 -46
rect 6349 -133 6394 -65
rect 6797 3 6836 114
rect 7311 3 7330 24
rect 7605 3 7624 24
rect 7337 -65 7604 -46
rect 7440 -133 7485 -65
rect 3831 -223 4315 -134
rect 4985 -222 5457 -133
rect 4044 -310 4089 -223
rect 3941 -329 4210 -310
rect 3917 -391 3942 -372
rect 4207 -391 4230 -372
rect 4281 -1234 4315 -223
rect 5198 -309 5243 -222
rect 5095 -328 5364 -309
rect 5071 -390 5096 -371
rect 5361 -390 5384 -371
rect 4280 -1237 4315 -1234
rect 4279 -1240 4315 -1237
rect 4278 -1241 4315 -1240
rect 4278 -1243 4316 -1241
rect 4276 -1244 4316 -1243
rect 4276 -1245 4317 -1244
rect 4273 -1247 4317 -1245
rect 5423 -1246 5457 -222
rect 6130 -222 6612 -133
rect 6844 -221 7706 -133
rect 7227 -222 7706 -221
rect 6130 -223 6153 -222
rect 6349 -309 6394 -222
rect 6246 -328 6515 -309
rect 6222 -390 6247 -371
rect 6512 -390 6535 -371
rect 6578 -1231 6612 -222
rect 7440 -309 7485 -222
rect 7337 -328 7606 -309
rect 7313 -390 7338 -371
rect 7603 -390 7626 -371
rect 6578 -1233 6614 -1231
rect 6576 -1235 6618 -1233
rect 6573 -1238 6618 -1235
rect 6571 -1240 6620 -1238
rect 6570 -1241 6620 -1240
rect 6568 -1242 6620 -1241
rect 7683 -1242 7706 -222
rect 6568 -1243 6622 -1242
rect 6565 -1244 6622 -1243
rect 6565 -1246 6624 -1244
rect 7679 -1246 7710 -1242
rect 4273 -1248 4319 -1247
rect 4271 -1250 4319 -1248
rect 5420 -1249 5460 -1246
rect 6563 -1248 6626 -1246
rect 6562 -1249 6628 -1248
rect 4268 -1253 4319 -1250
rect 5418 -1251 5462 -1249
rect 6560 -1251 6628 -1249
rect 7676 -1250 7713 -1246
rect 5415 -1254 5465 -1251
rect 5413 -1256 5467 -1254
rect 6557 -1256 6628 -1251
rect 7672 -1254 7717 -1250
rect 5410 -1259 5470 -1256
rect 7669 -1258 7720 -1254
rect 7665 -1262 7724 -1258
<< m2contact >>
rect 4013 3850 4138 3893
rect 5176 3850 5301 3893
rect 6334 3850 6459 3893
rect 7524 3850 7649 3893
rect 4390 3444 4431 3459
rect 4013 3393 4138 3436
rect 4390 3360 4431 3375
rect 5172 3393 5296 3436
rect 3027 2620 3070 2745
rect 3484 2575 3510 2783
rect 4390 2790 4431 2798
rect 4268 2635 4273 2640
rect 4315 2635 4320 2640
rect 4317 2624 4322 2629
rect 4351 2624 4356 2629
rect 7303 3593 7324 3682
rect 6798 3441 6829 3451
rect 6321 3393 6445 3436
rect 7534 3394 7660 3436
rect 6798 3365 6829 3377
rect 6449 2811 6490 2819
rect 6327 2656 6332 2661
rect 6374 2656 6379 2661
rect 6376 2645 6381 2650
rect 6410 2645 6415 2650
rect 7932 2528 7958 2736
rect 8372 2580 8415 2705
rect 3026 1726 3069 1851
rect 3483 1654 3509 1844
rect 7932 1729 7958 1919
rect 8372 1721 8419 1846
rect 3026 787 3069 912
rect 4824 1041 4829 1046
rect 3483 743 3509 951
rect 4858 1041 4863 1046
rect 4860 1030 4865 1035
rect 4907 1030 4912 1035
rect 4749 872 4790 880
rect 6873 1013 6878 1018
rect 4749 108 4790 121
rect 3937 23 4063 85
rect 4749 -4 4790 10
rect 5152 24 5276 86
rect 6907 1013 6912 1018
rect 6909 1002 6914 1007
rect 6956 1002 6961 1007
rect 6798 844 6839 852
rect 7931 696 7957 904
rect 8371 739 8420 864
rect 6797 114 6836 134
rect 6301 24 6425 86
rect 7459 24 7584 86
rect 6797 -10 6836 3
rect 3987 -434 4112 -391
rect 5158 -433 5283 -390
rect 6821 -221 6844 -133
rect 6309 -433 6434 -390
rect 7408 -433 7533 -390
<< pnm12contact >>
rect 6607 2488 6642 2496
rect 4548 2467 4583 2475
rect 4597 1195 4632 1203
rect 6646 1167 6681 1175
<< metal2 >>
rect 6445 5202 6453 5205
rect 3008 3893 8433 3911
rect 3008 3855 4013 3893
rect 3008 2745 3064 3855
rect 4138 3855 5176 3893
rect 4390 3459 4431 3855
rect 5301 3855 6334 3893
rect 6459 3855 7524 3893
rect 6798 3451 6829 3855
rect 7649 3855 8433 3893
rect 3486 3436 3886 3438
rect 7277 3436 7303 3682
rect 3486 3435 4013 3436
rect 3482 3393 4013 3435
rect 4138 3393 4745 3436
rect 3482 3388 4745 3393
rect 3483 3385 4745 3388
rect 4760 3393 5172 3436
rect 5296 3393 6321 3436
rect 6445 3394 7534 3436
rect 7660 3394 7958 3436
rect 6445 3393 7958 3394
rect 4760 3386 7958 3393
rect 4760 3385 5057 3386
rect 6206 3385 7958 3386
rect 3483 3022 3530 3385
rect 6206 3384 7785 3385
rect 6720 3383 7265 3384
rect 3483 2783 3531 3022
rect 4390 2798 4431 3360
rect 6798 3205 6829 3365
rect 6449 3174 6829 3205
rect 6449 2819 6490 3174
rect 3008 2620 3027 2745
rect 3483 2673 3484 2783
rect 3008 1851 3064 2620
rect 3510 2575 3531 2783
rect 7911 2736 7958 3385
rect 6332 2656 6374 2661
rect 6381 2645 6410 2650
rect 4273 2635 4315 2640
rect 4322 2624 4351 2629
rect 3484 2461 3531 2575
rect 7911 2528 7932 2736
rect 8377 2705 8433 3855
rect 13770 3510 13788 3581
rect 8415 2580 8433 2705
rect 6607 2484 6642 2488
rect 7911 2484 7958 2528
rect 6607 2468 7958 2484
rect 4548 2461 4583 2467
rect 3484 2440 4583 2461
rect 3484 2319 3531 2440
rect 3483 1962 3531 2319
rect 3008 1726 3026 1851
rect 3483 1844 3530 1962
rect 3008 1603 3064 1726
rect 3006 1500 3064 1603
rect 3008 912 3064 1500
rect 3509 1654 3530 1844
rect 3483 1230 3530 1654
rect 7911 1919 7958 2468
rect 7911 1729 7932 1919
rect 8377 2379 8433 2580
rect 8377 1846 8432 2379
rect 7911 1294 7958 1729
rect 8419 1721 8432 1846
rect 3483 1211 4632 1230
rect 3483 951 3530 1211
rect 4597 1203 4632 1211
rect 7911 1192 7958 1266
rect 6646 1177 7958 1192
rect 6646 1175 6681 1177
rect 4829 1041 4858 1046
rect 4865 1030 4907 1035
rect 6878 1013 6907 1018
rect 6914 1002 6956 1007
rect 3008 787 3026 912
rect 3008 -396 3064 787
rect 3509 743 3530 951
rect 7911 904 7958 1177
rect 3483 95 3530 743
rect 4749 121 4790 872
rect 6798 738 6839 844
rect 6797 670 6839 738
rect 7911 696 7931 904
rect 7957 812 7958 904
rect 8377 864 8432 1721
rect 7957 696 7958 806
rect 8420 739 8432 864
rect 6797 134 6836 670
rect 3483 94 3691 95
rect 3812 94 5391 95
rect 7911 94 7958 696
rect 3483 93 5391 94
rect 6540 93 7958 94
rect 3483 86 7958 93
rect 3483 85 5152 86
rect 3483 25 3937 85
rect 3483 24 3691 25
rect 4063 26 5152 85
rect 4063 25 4340 26
rect 4863 25 5152 26
rect 5276 24 6301 86
rect 6425 24 7459 86
rect 7584 24 7958 86
rect 3008 -434 3987 -396
rect 4749 -396 4790 -4
rect 6797 -133 6836 -10
rect 6797 -221 6821 -133
rect 4112 -433 5158 -396
rect 5283 -433 6309 -396
rect 6797 -396 6836 -221
rect 6434 -433 7408 -396
rect 8377 -396 8432 739
rect 7533 -433 8432 -396
rect 4112 -434 8432 -433
rect 3008 -452 8432 -434
rect 4281 -453 4315 -452
<< m3contact >>
rect 6432 5177 6464 5202
<< pad >>
rect 3740 4503 4296 5208
rect 4984 4518 5583 5208
rect 6170 4503 6726 5205
rect 7374 4509 7969 5199
rect 1681 2376 2370 2963
rect 9067 2308 9769 2864
rect 1678 1500 2368 2095
rect 9073 1478 9763 2073
rect 1672 615 2374 1171
rect 9071 516 9760 1103
rect 3763 -1958 4319 -1253
rect 4887 -1949 5486 -1259
rect 6072 -1958 6628 -1256
rect 7139 -1952 7734 -1262
<< labels >>
rlabel metal1 4379 2628 4379 2628 1 out
rlabel polycontact 4243 2609 4243 2609 2 in2
rlabel polycontact 4243 2625 4243 2625 3 in1
rlabel metal1 4409 2782 4409 2782 1 VDD
rlabel metal1 4564 2479 4564 2479 1 VSS
rlabel metal1 4265 2637 4265 2637 1 1
rlabel metal1 4333 2639 4333 2639 1 2
rlabel metal1 4303 2629 4303 2629 1 3
rlabel metal1 4353 2622 4353 2622 1 4
rlabel metal1 4411 2628 4411 2628 1 out
rlabel metal1 4436 2628 4436 2628 1 out
rlabel metal1 4513 2628 4513 2628 1 out
rlabel metal1 4692 2628 4692 2628 1 out
rlabel metal1 6572 2649 6572 2649 1 out
rlabel metal1 6495 2649 6495 2649 1 out
rlabel metal1 6470 2649 6470 2649 1 out
rlabel metal1 6412 2643 6412 2643 1 4
rlabel metal1 6362 2650 6362 2650 1 3
rlabel metal1 6392 2660 6392 2660 1 2
rlabel metal1 6324 2658 6324 2658 1 1
rlabel metal1 6623 2500 6623 2500 1 VSS
rlabel metal1 6468 2803 6468 2803 1 VDD
rlabel metal1 6438 2649 6438 2649 1 out
rlabel pad 2366 2389 2366 2389 1 in1
rlabel polycontact 6303 2646 6303 2646 1 in1b
rlabel polycontact 6303 2630 6303 2630 1 in2b
rlabel pad 6723 4505 6723 4505 1 in1b
rlabel pad 4986 4520 4986 4520 1 in2b
rlabel pad 7967 4511 7967 4511 1 VSS
rlabel pad 3744 4506 3744 4506 1 out
rlabel metal1 6751 2649 6751 2649 1 outb
rlabel pad 9072 2312 9072 2312 1 outb
rlabel pad 2366 1503 2366 1503 1 in2
rlabel metal1 6850 1014 6850 1014 5 out
rlabel metal1 6820 860 6820 860 5 VDD
rlabel metal1 6665 1163 6665 1163 5 VSS
rlabel metal1 6964 1005 6964 1005 5 1
rlabel metal1 6896 1003 6896 1003 5 2
rlabel metal1 6926 1013 6926 1013 5 3
rlabel metal1 6876 1020 6876 1020 5 4
rlabel metal1 6818 1014 6818 1014 5 out
rlabel metal1 6793 1014 6793 1014 5 out
rlabel metal1 6716 1014 6716 1014 5 out
rlabel metal1 4801 1042 4801 1042 5 out
rlabel metal1 4771 888 4771 888 5 VDD
rlabel metal1 4616 1191 4616 1191 5 VSS
rlabel metal1 4915 1033 4915 1033 5 1
rlabel metal1 4847 1031 4847 1031 5 2
rlabel metal1 4877 1041 4877 1041 5 3
rlabel metal1 4827 1048 4827 1048 5 4
rlabel metal1 4769 1042 4769 1042 5 out
rlabel metal1 4744 1042 4744 1042 5 out
rlabel metal1 4667 1042 4667 1042 5 out
rlabel polycontact 6985 1017 6985 1017 1 in1c
rlabel polycontact 6985 1033 6985 1033 1 in2c
rlabel pad 7730 -1265 7730 -1265 1 VDD
rlabel pad 9076 2070 9076 2070 1 in2c
rlabel pad 9077 520 9077 520 1 in1c
rlabel metal1 6537 1013 6537 1013 1 outc
rlabel pad 6625 -1258 6625 -1258 1 outc
rlabel metal1 4488 1041 4488 1041 1 outd
rlabel polycontact 4937 1045 4937 1045 1 in1d
rlabel polycontact 4937 1061 4937 1061 1 in2d
rlabel pad 2372 1169 2372 1169 1 outd
rlabel pad 5481 -1261 5481 -1261 1 in2d
rlabel pad 4316 -1255 4316 -1255 1 in1d
<< end >>
